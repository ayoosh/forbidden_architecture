XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�<��O׃E�︽J�b)�������^)u��;����+ˠ��[EuZgfĜ�����h�a�d���Oz�P��O0���\9UL��g���E���Q�en_z��YcS%y�$�a�be0�i�ƶDKG��ٮ�hT3+B��'!�.ۭq�i�ix�@� �Ux��E6����iK�"�!:�y�#�`C�i��x�A^�����5�g��P���x�����cT�3'ڐ�oCj�
*x�٩�A�fڢw���3����B������v�X+�Ĩ�]�p�����r�ɣVN��,�=��!�ޥ�8�uU��N�T��X�|�*`ռa!<� s�y�K���K�\�^��Ƭ,4�sN�}�q���ҧ��ے-�		-�w���f�O��Q5�n-̘7�9*2��dZ
񸡋�n�u �\�E�G�
�b��4>uZoX
!��}\R<����)Ykl����@C���QＯ�aP��i�}���󷱹ʑ�>iO��]�6O�e�"��A'�x����>3-m�t?��4��+߆�v�p���J�Y����7�*ǵ�-tq�2҇L��9 ��/r��8#����[zW�#���L��o'nqb�އo �����,�Y�|�͐�#Zi���?NI��������D$�q23{u��~�n�ѱi�� ���i?�y��������e��!�/8�=�دeu�*p^��"�͞C�OU�^L�>��B����S�lK}��D�d[��m��S�t1XlxVHYEB    fa00    28e0��8��*�¿�?*K>���:���dP��Lm�72
�T�|瞱</�-���
��l'��6S��
��@2�_0�Vw�Q�AR�������R���y��o@e�J�� t���yq�w�
>�.&������ۗ���,���D$+lp�Go�Q����\�����un�01~!`(��:�Ue�ܦ��\����KS9��n�Y�B57u�8�Z����Ï|�H�ڎ��ʵ����L����HD&(-����Y}�(��!���ۃi��E~:1����z��%T��ĕHe��>k��ɝ�X��@��jh�{^Θ_B�uE-�~��ؠ����ˀ��_�������짛c��e������
��'��̩k�֌�ȥ+4�@	Yw�W�WR ���9�жB�}�<{�H?G76������9�=�B��B�?��5�!�fe2�xS�%�����1։�ίJ������[�;�*e؟��#HH�%��^�`X�j/��ɩT�䏊gP��RA�Ĕ�D��r#c��0�2��d���,<o^��#�|eڤ32E���yk���ݱ��%L��ㆻ����[�P
�Q=���\$u�NA�}p-���8J(�3o��cO��R��O�ly'��V�d2z���K��"�W
L��c�-�#���w����QY�J&�g�kI�x��mby�2�{#Qh��_v�Mŷa¸WB��zw�jY���B�42g��A�	[cȐ�q�/>��2D����bM�H��V�O����s6i��Q�U�=�9m,�>3�Z=��p���ܴ��<2��}���7��}��ĳ���R�h��C�ɢDG(6��-�v�VX�K �}�����_�N����g��@ES�b���ጪ���b�]���Mi��_䠓��_����l�N]�	4'ZڛuRl��Y�\|1,_��8�[)U��d���:c�������*�oGy8R�gL��$��el# s���z؅pnn��fe�����A�3@��%:�M	`O�k��p�L)��J�������LΖZ�FNZ��u��Em.y`��[[�u�_S/<K>�A���v'H�co�S�j�>$� ���**$1�ͬ_XOa�*y?Eԋ�]u���-�tc�W�@��
#�pCmM�WR��j��'ק���.)E�ϭ=ӑYq�P�

w�u�⪍���O^�/,~�5Qq�"K�-!�Jl��)�h�)K�R^���3n�&ٌ��=���|�l��n�i%���*|p�5�v~��7���w���x�� B�w->���~�ֈ���@S��C�H0�P���c'f�a��:��i�I=�S����,_�RK��������!��r׳��3>ҷ�ϻ��7̾�l����g�)cfq	ƒX�a� ���h���I��)�%e�+%>��9m��ҁ�+���s��l�&�ڝ���}�Ƃńlg:Qׯ��%�0tS�v�xѡK��:YO�q~�]�6*4/�`�4q����+�dh�����E\��\Ϗ�̼�&��Kp��>�H���](���GEB��WW�2T������דj0�A$Qs�}��"��rԭ|;&+��E,- �� L��B��	ȇ�Ϣo���������#����Y��.V~�Il�������A`��姇 ��S��}���I�e�m#Ġ�����)�� �[�M�}B͙�bQ�����b�$�Ꞧ�SD}��j��;і�q����dQ����B���TѶ�]�K�%Ҧ-S	h��3Ɉ�-;�o���+0��p{�F�uzi� u�}���6,;�j��-I�pUx���ϸ-I��Sr"�yEgŌ�L����^��a�VuF����;D}R{a���Py���=~[Q�e��PE�������&�_��pK]4���Exx�Ā�.�n\�Q����z�ߙ�C�D� ����I�G��:$1��md\�Zڛ	������︓��B�&U��^R��x��1>��C��?p)�O��CG�N�4��e]�Y������iG����,�o��nm�������N��'j�ZB��K-ӭp�R
`���M"A��Q7X���P��=�L{��:'��F�r h��V�Y��# <�>lO��YA�Fl���DmQ���;V3�)@��$�=?΁��ue���pd΂�BA�Ԏ��x��2�b��]�����6�JٸY��_mA�	�	�h��=PO4���7�"����\[�)�s����Vl��E!.�a��R#��(��>�1ot{�����|ᗢ-�>?v�e`����>qGO���.JF�Ey�@��s�.IC�ty��O�ʠ����H&����"��JmH�,�Ŋr�pm��3񖦳�o�{4�{����[V�|fp�O+s��K�8����9Px92Y	n~-:�DI���)g���baU)?���/��h��C�S�H�]���)Zs�gz��]5Ȓ��{.=V\vl����b� �ʍ:`�b��ǃ�dj��N��:�P�$� �2 �I�PNN#�.�y��j�m�;�萦�kV/Xn��-�M�b6$����y��{�+~�tx�d���M�:�=����Z��Bܱ����ȼN))��d�b=���~[��cp�t�&]hcfC/Y�2�s8)!�{<��CU�� '&�(�I�\J��&���*���:��T���;�N������>g�	�u����oXy�섋�9Z he(D�M+��Q�X��ɇt=����e�wӖa�=�IQȎ��ׂx<��
��}C��9;�iL���rG�e(��SrR�%�~#�0�3�k��|�]w��w�?E�>��u~mcaw����C�!\�Z�r�ST��L��|�^�@���,�q_�������B6����DF��3�ӂ=aw�X�O;,�	!�tO,�?v>���N���`D�#��#�Oi�6 QĽ��I�3�2���P�2]�&X%�_��G����
��� ��f5�<spB�����#�ș|����:C��T���J%�w�a�)v�/m������@�X��X��j9��T,ˡA�%�C�x�w����zQ+�\
�j)�K�3���ʢ����
�0tE(̩`�1�N�%,��X��3�=$�0�kzx't��Nt�Q�"�	-d�\Ix�ol�~Y{>��:}��3�*���wzZo�F�,!���85L�\R۞T���_�m�������1����ւ�s�L���6巖/&�ρ��\���F�jV�
�'G�U\�Qd�6}���T.�4[o��?�uE�:��$����\�"��gz�c��p�ѓ����^h��>S�C��M��~\��FTxb���q�1�s6�Qy,�����VٝP��h���➮�O�C�D I+b��%�t��K^���b��Qx8jG�ZM�i��ԾZ�9`,-R:а7�/i� ����\�_��͘D��M=��n�
E,����� .߂�N�~ki:M{�S�Wt"����U���ۃ����v�ٗ��ĺ��v"�K�}�}wT�6?N4B t��f����G�3�Lգ�id{nҠ�6`}q?RI�,%�Hz�*��]N$_�g@�D�����t���Y6&4�h7J��u�RЕ��*8����5���j����%�B�̮�:8t��i=4.[9�"����	�6Y���$٨R&7�t�l�(=m`9�����E�h�E72v+�l�K6�,���hȒ����@&\p0�r^Lٜ�7�i//^�͌:m����	���<Syb?K��Z�u��R5�ϻl�z�x�1���)�0��L��ȢQd݂̲��+�"��d�r��F�aT�Md-�u�7�^�
q�9�f�0&�����q�ɸ�/źT �`'�&�"�n/n�z�N\w�
 ﯗ�|�@P�����,��}����_FH'z��F#�p���l��5�l�$���t���{-\�D���2��>Kf(5�HBz����˪�v�3�:�jV����K7�-���Y����8��zh���S�����jW%uL��喓��ja�(�Xe����E`���bJ��L�~��b6���o_�H�}�[]]��ZhmAᆜ�:�B5�h�n�� ��*NG�_�`��g[��$���!�)�-U�W�<蚤�~�8	�\�޿T\����vt��c��� 8k���{��~>K�Ŧ#�S�
n���y����g���qT`{	�P��~�cf�>G�P4!�!Ry)gkr�y�� n@�_�f��=���9]I�1:#�,H&���ӷ�����s(�j��A�!g���@�2;�=*�6J :�jZ�3���}�[u�&�/�?e���ޙ�����ϳ�y��'���df$1������N�ҽb�||��{	���x ��h���'S��0�� ��`!@�?pjq�)�-����jݖ?5�>�-7�@b�E_K��������'8�f��2��z��&�xxL~и����s��a���ޮVC����Z�1^�T;�	�^�) qIpI1:lblb�L9�`�L"rڲ�,�Ԡ��Lw���QO�}{��Ҟ6��A�o�"�[�a ��=X��/>�+�Zu=�mu����⁫��� �jkuGq�H+hi=!Y��nD��ߚ�M(�-���w�괾v�!7\փx���X��c9.ab�v$0�eW��&¦ A����:�c�ls�v�V�JM]K�%
g7%�q��J�D��'�$�ײ�,.�*�W��lD�!�P�K,�bG�>��G���c�[��
F�g��v�ϑ9��@w믒�4-�$5���q�2�
ٜ���h`�$�I�)��2�P>O��ALD���*dt���V��/�XT�<p�����L� 4,��G�dN�)0g�z�S��Rm�/f�=^s�����b����r�G�b�N������/HB�>9�k���例Yδ�������+�ɛ����C�Fԏ�}N�H�Kp�B��?Y��J���r�bʣ�d�_&Pf�9��QN�Y����[�6&x�LY�5�o����w|�F���<+&�9�?,EN)��ʍ�cvK��x���VO-y�������ŘF$�� �]&(ά0��]�jRB��*��y��S�$�zE�W�u�H��e*gJX����X_q��j�8qh;gr3�Ҧ�[#3s&���Љ3<�q�2v�\�!/����\	b��n-��b���
G�s�v���yڞu	�i@qnpeP��7i��x�н/U�����_�T��ۖ�"�uA�=���� ;DƧNN{Z$(�Ci��2B������7�J�Hӛ�f�B
��L��?9w��/EI�K"�t���*��p�F��ok��`�,O�{�.R�%B1�B�0X3��r��͖��&��א7=�?k��_��TH���uJp�dO�ќ��>*I��v���&A�A�֕8������[���U�`��]u���aF���ٕv���b��n1���s5��9���Ɲ��fo�*����S�:!��Q�\�Z3��~���7�����$�^!i?��\!�HՏ�GՃ|����\�5[f9�t��	�,� D�&Ъ�&�
_vy??H�����|�>e�V��>OQ�Z�+�|v�����$���+���ů��V�W���?b�=�7d��~��Ư�+ytQ�����q��Q���Y-[*lpBl�S�Q�_,����Yk&���a��c�{�&�H��j4f|Em�z�:��1��>�=?)��Q�V�	�ZZ���Ռ�ߞb�*`jH#4X�.�?V�o�� I4��=���n[�x���F:0��&��*D� 0n&�x�)�>��b/�vUzWi�?�q������@�M�g#
��GFњ��4�}��' ��I��)�u���7��!�+�8QOtP�0���52�r(��MwmAZ��uF�C��6M�]Ebh*|���v|	`�"��0�����-s
�	L�+g̀���K>��<y�r&�P��F.|r�\v8}ݽN@�U���+��UQGt�_n�R�:�7�*����eҥVFX�I?~zt��1c�o�����^�`y-F����QS=�5�S��="�J�L����T�q>�CD�f�{C1�p�2�urѝ����$=Na��9�|�q'��>k&}hu��<�~.tA�1�0������X;X���4]��#>&ա�K�ľ|%��@��.�_ �0ⱍ�{�`1}� E�h�&�����g�ů�/:f\\%����|��Ǆԅ����[�C�H�{�۩oR����"݉ƪ���B&Ҍ8|D�鹶0Y�5��+L���֕�^f.�C;���-��E�?ٟ����Ȳ� Y�֮g
�)�4xw}%L0MÈuz;{������Ir̓{ �����՞����A���&�KYpN��t4������r�w;�!ħ������t ��X����w��0�B����#�a��Y�9������G��[A)Z"���O#����Wf�H��+����&)-��j��00��+�����R�,�dl�V�� T�J]��_�)�+�J�����T%��駢�J�B-y�U<�ܮ�O챑G��¼6shz�ڳ��)�Ղ�n�1#�P�@f�%o�sJ�;EFakk_�+����@I-ѵTR�cĭ����z �P,}>ye.�	���5����,i�,�R͵!c�^��3��.����j�����Qs�A��-�lS�)�N%�m=�,P�䡻n�t�5�Z��$�FQݿd�dEz�/������3ar>d�E�K
��$r����`��O�a�Ax7�x8�u|4/\9
	7�#�r����e�i"�t�a8�6��4�x)��/z������ח'bi�;ʭ���˝eqG`��Z\0��:��˛�3�Xf"�+�l��,�E`5*#�Y�i=~�:��� @y&� ���]�@���ˏ(p�#�N�lfթ�y�@U�q;���%�� ���R���D��"�ML,��Z\6R�h���x]
_E�;ĪR�ď𦮘�����e-�Z�,ϥ���k_���f�!��xa�ac�����ʻ�>*у!����R"oS]]fYa�ؖ���V�|��/Lk�7M�ރޚ��/	�M�ͱ)!Q`�/W��%�����b�����D!�hu�����]#T(��# 8(�h����W��m��5����[�^A]�Y���zy����K�P�6�B�pvD��Q�����
�2kZvJ�?0�4P�B���]̬�w?�΢l��&V[^��\܆k���"�ŝ�B�V���yg9H�N<e��������!���m<����� �Q��t��Tiu��α<}�;\�0E��H|����g��.ܬ6TL�d��KЬQ8��&�ɒ�t�Q���/Qݭ;��� �7�P��	-{4n�B���˛��D������	�gJ�6%aS���~@֏���s�H�r���ջ=x��>���5�H��sn�B�a�FH)&D�0+�WB+O����hQ;8��Rb�Q�G^�l�G�S�Ţ���K��u{�4@���u���%ۮ�OЈl��ls���|n"*<��Fn�%';����0E���`�u�A��4p9�L��	8��*�6F��_��nW��s�)��kK	��Z������u��3+��Z�u7���f�<��@?�G9�5[|��S	�:�N_�N-o�~�?�6W¤[uR$�,W��C|�Wy����^�f��6�R�2�����q2i6�u"�S��<nYczH�M����b��D'�A�Uͱ���V���F�$HvĐ$]��4z9�gf�]�h�R���;wQڊ	#���((�~B�u���Y"a{�G%2��+P#	��S&�bN>��:[1r��N?���"	,G�#���~����9���,��s�1�2 �p`Jb��:_?zkaY	�I*:+t�f�2+�a�A�\���Y}ʃEb�7�@A�������4ځ���4Ӄ�;g�w855e{���pn�Gy���[���+����}������̩��VC���g�ٞ�?u�a����eٕ@��l۟�"u*��y��0׭~��� ?%��O�yE{���+ܫ��o�2^s��q�D7���P6�Qj4+�8��Pn��}q3�0H7�|��qK�[#Wf�{�	a�2<�;�7�J�{������0�j󋵰�/uWQx��pZ088m����ޙ_V2��.�5ц[�����u��!o �B��v�W�:���uM�s��@�h^M��=�-���~P����%��k=[����V+�ݭn�7��	����|:3� ?s�$����+��y���v��Ǻ�`4ܰ+�sR���͜3$�X�ʐ� o�y�S^p� �xƎ���H���|c[3 	Ū܌/�A>�<F�BkF�w@W�D�ۮ�����(����㎁�x���BHуp��\0Ne�i�@�On���F�0��U4CmR�wD���;^Ԙ��2�XD+��8ǘ@�|i-vA��� �?���$���s1�_��Q1��ք���v�u��
��kKL�� �c�׵n��I/rW���*}���3��'��a�.�!̓�r=�>K��OZ�L�p�r���(�
<���_�c��iúv�T���+�WKIJm+��|��b��~��0�B���ݳҁ^�G�C$��]H?�Vo��1,�M��ٔ�J+�����X��иOg�����W�C�bJٍ���&��� ������t����2�N�͎�*�Q���]DE�=mƱL����,D"�-PJ]T��F��.�;o��e����xPPPHc�SSd*�10��7,��S{>E���qF{�\��� O�e*�l$��8ǘvV�uLټ�K�7tNh�%d?�W,��u�[�ŏy���u��pT��/Y]e����h3c�.�ᒶ,�5���_C��M%2���V�Ӛ��x�:�!\ukd��SV��D�����3Ki�����qj�����bK�Z����xW'���c��x�=)��g*+�T�f����N�#(�w���ʅ������|+�Y��(�R~�X��"�Tyd� �L`��ǫ(R�: ���zj��x:UQ���R�
܇C2]�t��� 5Wx���Ƿ�)1�~�Eu�p3$ç�8��?���,���F��*n쓈saNgP��=<{��ܺ�yb�#3Q��R:`�"�|��rg����,d�vK���d�o{�^�2g꘷
�f���,���4�_�2G��g���J�x ���_T{0��Xά�Ƽ-d �ո_#R�w�]3�;��o�c�\��ʨ�T�b�aH>��N�����9��2�UG�mЋ��<�=]'�˯��]���_�Ow��׾vY�����)����\&X�R�x����K�'���(Oշ
:�Һ�:�	y����G��)Vj1h(P&k�40)� ���s\M��#��{�1���b9�?�*Ҧ�?�8!7��8*���-��^���Y�?ŏhڡ1"�g��G�E���ٴ����PL]w��A9#H>C�۔+G"�2kf j���Y{���ΕX��s�D_�ѥ	P��S��+tJ�B�_ő*8i����
!�긬�ۉ�@����@��bH���Z�u���G����%4������V����`G�M撑��k�y+��
� ������1h".2���S݁n��uA�Fea�N��n:!�A����{�F#�ҽ�B����|�uC��%r���!)�{���xq��-��k� b1�=IU���a6�j)��.��ƨ�Ø�W��WHv~=Myb���
��?�fA����/g��'v��\�(-U�M!�VLd��Of��kV�����WD�X�L�@�f��e2��jVԟll>O.�|�;�h$<#L�Ýi��85��&�;ܱ��h=^���N���������K�h" �&��j�vG�ʡ�ߑ��^��2&�dȥs�o�p�4��>.c4]�����>�%�:�>��N�+���I��	9+��s(M��("���kn��(F/�!T@,8V+���ڰ�n�!	&�B!g��q�xxY���x�q ���e�a�l����R��wuPؓW��o�ߋFt�69K�D������e� jO&����{^�Z��s�Zx���n�>5��~/{�Y�%�N���c�ca!q�sL�o��PoN��.�Hˆ�ٷ)��='��bZ��w��1H]� �~�K|[0�kO���������
�٪n���R�����H��G}�T�@�J���X9�)�8<�����?�Ћ/��L�ѺR�#�s�7'��XlxVHYEB    fa00    1d804mC��5c�Zr)tR� Y��� nI%�����v��^�'�w'� [�PU5^7A��5zD����06���H����g������A��u��&��L�2��t0�8s�A�c��*YO\�4�8>{*� �Y(x�M���1x�W!;KX������~Y)���]A��x�5���^��wD��o�������Г0y�_�����v�O�ݞ�U0%�c�ް3m E��+���G�Y[l�\fqq����H�q�0#bv%c,�����q�&;���������j.��퀏���u?
��,+��8"v��������i��^7��~����6�%�*�,z�TV�*kƤ[Q����)%{�~�"V���	�;;�|xY[����?�Xrb�Yr�8j������ĥ��H�]X���WG�����_�~���,~���ѹ�\�Ul�R+��x�q�<�J	�',V3�\�r+R Z�����5Q(l�i��f!V��s�0nu����в�R��r\����2�2v-��O������v7BIf�CIz"��M[���挝��>����.�%��sks��|>�i��F�e/E(;�w���D�&Z�hǊ��?4Km����[Q+���u�1�Ѭ���O3�4(8�H?{����Ah�D�Q���͖l1�'��_Ȟ�,/����%l�������x��+�^�I�^�=IX���J>�+(�m�ER�9�� <|?�j{l�%��e.F�vҾ
g�;����T��l͕6�-OѤ����M�;�%*��J��9�T����|�f�c
56n�MT�=��f9�~�X����,��N��k�5�kEө�R�1`#�Y�К2� W�ݧ,^ď���!*��)�����4	�'ѫ�[μ�6��)�����T��ƠӮ,[��$%7���a��?��ͷSKb=���.�:JV��o+��$�M��&8���|8\�l1NA%�m�m�v��:���^����菖�ޢ��8u�K�/cհ(�x��zZ�@eޘ!��[�A-����e����6p���¼�"�7FUh���Ws�\��i��z���ŝ(	{�c7��0�sp@�� |y��R?"�d���.?P�`h�Q�E��3<��t��H���o��O�
U�G���N=@�U��H��WŬ�l������GM�am$���_�+�o�����:�+_�I����#�Q�OP��L������#��;A����2���rQ�1"A6��tov�9H��-�s��#A(c+W��hżl�/&�h��t���~�.���\f^U�o0�qrV�s������	��(h��xh.���4,jV�����&ɧ�Z����S��C��*u�d�O�����؟�Kɵ%�d]/��J��vr5�W48�0u�����������ƃ����t�,s�����%?���ۻ��2z���oE�Y\�韾/IR��W�Bh��SXĪ�j�J�#3(�B:�'	5O��[�ym(�u�S�Q_�W`���w¯*�?�H4򘰉ʴ����f�-B�~O�i|�i���݀V����b<\���Θ�'~����J<��� �1SqP	ʭh+���3aw���Xp�F�Z��-�
N�½���u!��׾�-���Pc�AP�x$M`̎#c\�ٯHp�E��=	��H���_�:�EZ�]..��?GR�=j�̩��(��WK�!��~X�HUc1{w��IF�n��>�0K�,�v���;��7�O�� ��#��!�pw;7���wW���v)��6϶� H�_ _5�:Dג5�)}ܑ�H5k�����~~�Q{�j�z�Q�;��"�u�u��_`t���eU[���%+�q5.Y9�e�潘86�7�"��A<�� H@���@;E$� �Y����-�>�Y*(*
xB�1�����ώv�=��C7�N� �;��i?4)?F�_	��H�,,a��72�j���A�@4r���a��4�X��4��d�8�g�� ����w���"F�*���'4x���$N���;�����n�+�u!�Yf;��;�шK��>�E��.�rqk��.�#��Uq[��=�M���tf*��0���}��o���bC�C��L�Y0��
V^�^�E�tM�����Q�\���Y���J4Cm9±�$��Pu��{n��n؟ƺ�U�P�_g>�@��zR�;�M K�FY�ݼ�]SLÈ�uZ�G�Ǫ��3 0��AV&�H���O#&��ڑ����h��!�O;'e�
>��{��p�3��>�����.U��MQ �t��
�u�1�Y��-�ۀ�����{�;@B��W3���~P�|-�����9�$��"�i��_�bxS��8��zL��J�%�>q
6V���Z��b��~�~i��'�C��D,&Ey\��}�3S�~
7�F�OITLkm���"��2�i�'��
i�:��Z��1`WoWs3$�Y�.$�-��jo	Xiw�c8��(=�ѫ��fOt��q����U��c��J��)}�?����ӽa���+�ɲ��+F��Pq�Cr�Sc����q0B��+�D�.�\�[s'I�o��~)�:I�CI}5�քoq�g� �f��*�|b����ߵc+���ú��&��Jϊ0��J���T#��Y�/�e~�?�,k������l�J<l���=�(�"�����w�ތ0�����0��p
�u)��=��@�5���{�s�{-Cd�A�l�/�x�肌/��FH�_��:�s�5�<�-��;>
]��G�X�;�d`:FC(+�+�W`�#��Z�Qol)��R����]7��_���(Z�	K��<7HoUh;��	��)�8�n(A�˱m����4�Z9�%u� 3���/�Y]��v��͇��KN���"�r���n�UV��@AA���Lud�Z�nYO_������|j���1�)��{�Jp�T�ӔT�|B5��D?�D�^X7�rG?�~ô��i)�T>�PD�����ٰeM�mG�B�V��|}q̚	�B�ua��������G��ʒ��s-�|�.���Cb}6�t�u��f��f��c� �yiHa�*��	���C�QQ���;x���lx�?	�i�J���Pi�w��Ȑ8S6G���;"��?W1ŅO*�TL�����6_�a��YR�Q��b���8��;8��= [ʤTDn�={���+,Gk�cĿԨ���ҦY�<d������g�*�+D�� ��v%���'��y$m�<���dHC+�����jkp�JHN�l%p�La�^j3�Ӱ"s��$�ģ7����/HG��3����a��=�:�}i��K��'- /�Xg�[7QS�8�MA��������_Lvo��H�9�5Օ�p����lm�LDj��L�O�ǎ����=�`�F�ԑ0;�gK:�;�1�w��~jF�ʍ3f�pNECx:�W&�$��(=�?F�cDw�][�G��m������k���paA�-��H!,������BOVҡD0>MP��/��I����7�����g4��C�F���c��?`#s�&�#%Z�*4Z�p��,G4�Z2��Ov����Q�p��g ���?r����D���f�̣@<�z��5�$���N��=q7�n\1�^�RMUQ�4�ˀ���`���(��/� �K;S1�a4˷���%�����1 ����*� 7ނK�%��*�J<�_�� Cx��\s-C.���q����3w��Kx]A(@�gԲQ�vH �@�(^39~�����j�A7�H,�Jc���wY�Z58���!��݊�)ga����GSGE�c�����^�A󩂝k5����ۗ��r�R>}�l�f-;5�o���3��%'1��_!v�q��8���2N(�y�.1���7Ii�R�|�o҃w�DT+Z���1p،EC��8���xOw$b�b����bm��>��LCK���
�۱�h�����A����kFa�:6Q;�طbNE.Nh��*G.�el�B1/�W��b�abb
_���Q.2 ߡmi�|��:d�2������̑=�}���w	���>.n-5ϴ�N���BX�/��T�Lǿ���$�}\�LH�j�޲z<%0�lH�~�4��v��A���Ϣ����Z���m���#~�nݺ|��Ej��l���|�d�@e��D#���M�M���Ug��|��ӎ0�䥇֊}�F�K�ĵ3Dsk�:z"�v� u��*��_}���ߓw1�ޑ��I����<�H{�2���ݑgv��[swD�bO
���<��,�Ʌ-� ���~Xd|�i�>s���\���M�����-}%cK�VR(�����W�T#�핉pHyз�I�s��4w����v���:�<�y!�� }["��툔6��>j��)��UAZ{����s5Z�C>���S��I�+� 6��n��/ׄ���&�v��H��=y�[�ۿ�2h�����b�vp�wdrS�-����Hh4��✃�߁Q��(���~�������ʇ?1f��l]WB/��K.&�eW^� e/67��Z8�/�X���XN�C��}5�� <�J�{Y��T
�f���x�uΰ˄�p�׎�]�R����:�7a���z��l�΄��A�1�t����q ���d?��K� mEJ&����9�o�)>*��WC**���NMMZ�Zz�]dա��Ԙ��@���9�\mT�S-�+T)�r����܃;ضZ�3�A�����ps@3'D4��-��w��H�8�ڤJ/���G�H
��=�� �+�Bk��#.6.P�}h!Z���^�	t (����S�������:�B�g����j�R�l��UK#k�B_�?���OWd2�S���{~=պ场��/(�>i��J��X�TJ����t��Wxuy(�z>��?
ZC�0�&���r8\ET�ut~�`��H��,�<��/a84r9
dV��I����*��_�$���zl�_r	0�,��Ȗ���ך��}f2bwv����*���ؿ��/t�qL�m�,�S�� ��a�P�i�z�����QQ���>����O3�q.��[��yv�m�;jQR�xα��4\Y�&�<FU��&���A&��w(�W�K��Ŧ&�)6�����Q���k�:%��h��6���\���Tji^A8e1��6	7��(݃|��9+�}T�|�A$��t3u��� �q��.c���}�Y�r"���h641r���L�����Y��\�vsӲ�D�W����A�nY���9�Qt�����IN�'��޴؏(c����mɓ��@��o��Nj�5*����q�G�Ɛ���Cr5;fZז1̐C��~��q-u��b�>=\��U!Q��&���>�j��^$R_���~j��0���zQȌB]W����ĸ�Ф��TJ	��������qҔ�)�>_`%�M��i<ѻ��Y&����8Ք9^wNj���S��XO&J�����7n%��d��S�"Aߟ��� �%0r�O	�w�=NJ���P�D��W�v�\�\���/�.�n4�Zw@�N�6X�����`s��}v\��f�HJAɼOz`2��ƹ��I͐�3�
��0�rU}Y*d�O�2h/���h&	L-Dc��j:�df�Δ�!yh�{�!��e�:o�O������������Vv��_������v@L܎��%'ۉBTtlHO�w����҅hf��P�|�r�o ����w��Lu�m8h^���I�rB�B��P��Yڿ:�k��ȑ��a�q��sB�V��"�������	�C��`���G@�Jڏ����h���T�@Fw�h�:B�n�>g�K���	#���G���}�-c�˪�p0�+z�{�sQjCW�|���PA
�טxZ�ذ�����MoW���������y�&���~���%3�Ahn�����P�k����`�-�  ng��M}3���O5v7�>�04�pF�c�y۪Zo<?uH1��QIU����S�f��F�T�R���I���a�^!tiKU���Jج݂lw��'��*�m��uKN.cъ-0��]	��&�@SU��&�+�0Y�f���2$L݀&�M�i�д#~y��f�t�i��^���$1���Z�\}�Ȉ�sP1}��O� {H���9T�@M���;�tR"�"��g<�>#`y8�>��5\�Si}�e�_�&<�F_���(T�4'xL�����6Y�5Y��u��O�@G L���IB�Xlڙ��?��wq��I+��>�g�l}�TS�';�t0rgwB%�4ݡ�(b����Ȓhy4�r��c7�|��(�7�m��U�z [��}x�������v��u=�	{���'���l�E��X��+A����۸�r��C1�xL��<�iu���10o�*�d��/���$�`��tE���I����yv������`�� d�_ h7�J���R4v���w�]��Y���J�[������L� 8[��4�\����{D�m���&�LIݦ9�s�ދHM�a�7��4[�ݷV���w\:��E�zٟ~�%V�-�$�X
<h �g����5���^�8��,�2�Ǐf���P���;BY� �+���W���<�j��~c��vLj��J-VE&��QY���
��gQׯg]��_�Oغ)��l?�M��|������g��f7h����ܵ����>J����w���HB!����gqP�w{�����E쟛�-e1*��b�d��Ts��[(*�G�-P�
�����t)���"D�c{�vL���Zp�ˆ/��իrxk.^e,~Ѳ��z��c`�1ڔ��d�
�l��F�@:��UМ��)�I+�F<G�9�)q���ZR���U�hT@١�'���"|W#�͹2*L��x�5d@�·_�����Z?$���_��V�W�:O���������!�l��ɸ��z��:Q�k����J!+�/�ُ�3��B�*�D�I�4vph|_������J\��QT�R��<�AQd����S��Iw�A�{����)V{ps�h�es�r~��q�����`q�pBҹ�P%A�B�Z\d��wu�o��k�{D����*�9�<(��rݞ��hs�G��bIѓ�y��e��,F:_v7]��o�뺐�=�DDo'h���΋(B�*���1ݨz��2U\l�_�X��)��~����ܶmF�j�ɺtw�׶չ�m�zL�S�3�\�^&�sZ�LC�6$/�1X��d����jG�2���u!��1��oO!�a��L��ӽ7���s:ߦ;-u�UF�U)�7���w��R��ݐm�LGx�����NJ�e%�|�ʏ ����le.�J��s#�l�����Y�0��XlxVHYEB    fa00    1e20�uR�8�?���iQ"`C-:��5Fۜ0��+Ki���X�HM�����D2�5<� b�o�	˅� ��b⭓��B�H�����	�~��#Љ��`3؅��/v�/��3���,N�Ǧ��3���'{<5��Ƈ����;$���>A�<T`��$��b��Vٶy��{�E���_�v�*��,�2������G8������m��ad��ՍOU���|�߳��(��䶔ÌI{��N��n :�Lj�J�*��M$S�8a$Z\��sa{��@D�,j>j�v7n�ѩ�@rr
:��ѣ0�T�,T͠��x�����}��@��j��n5���%4���{�*�d[�熫�� Y���)}�[�<�>Vj%����Y'���A�R./���K;�[F%ڍ5D��9����,'�iZ�<`���|�n
���J�<
ء3e&2}� uɵ��o�yI|�a��bo�g��a<�s:)���m������Y��i^�1�*䷐�+N�yG�3AݧnB��Xxo��,�$��p������e������wl�KR��$���ky1�(���� ��:n�Z	ޮI�͌U����9x�p���r��TX���5�A=K��I��6N��:����m/���C��X�1��6"�����U�O��qx�5�V�3gzڅ����N�+�,G)��P%E��* -N�ȶEF� }�[*񦟐�[�&��`7���I��ֹ`^6�K�����*{G�K�?]�� ٦$8�U��j�P�Y̋��H�4���.�W<�<���,VD���"b�+��;f��m+�%P�����=��4Zf���Q/��s��?��9ϛ᫊I6}����vq�8�ь�
��+T�|j6>�AptS1�R��Q��d���E����p}��Ij#�4@��+�(I^�˥����]:�t��`H=
��5t��<�.�u�ͽ�$U��}�����;_�wWɡ��C�.�;��Γ�bɐ�{8��n6n�۳�/�5�LuX�[v��aH�n]�ۮ `�5G�.S��\��;B��7�OY�s���4j�{�Ng'�����,��q)�^���Z�Z ��jS��S=����[�ͺ�,�L�e�%����Nq���c6�݅=�k�5���l\�!�Y�P#�z�hf{�m��k���t�sr�b��O&A5�\�����Ѳ"bH�����'�+���U��wI�.�80ԋ���Y,�&������|���J�'��������q{��Ş-��P����CI���B�F�{��O����9Eva����Bx�8"�4�{9&���6���K�c��I��^�υ�҆{B�
uʚ�7Dd�	�G��:}H�ا��tG�{��g�V�����[�!gCQસ"=PM�a��oͥ��b���+��=�:������$6Q!M5nk��,���� 4���##̯�8a �
�7��y��Ld#(��G҉)�����k����c��.��FX��K,D��Z��2�6�NO/�_�1�F��5���6u5<yjV�ok�e���l䍸"hޟ_>���Zܬ�˓�N����+��H�vNH��7�RB�v^���ͩ�*���f���y��7#��y�f^ك�����j��P�io�i��Z�c����cY�J}k�m�R�JЖ˲m�K䥨�'�)�X����Ks^�<.Ϥ�?�ߠ���л��ޅ_pTG��a[]I=��6�w�7���F ��wt���.�Q�_�>�5hy��E�d��]�a��c��ܻw���F�C�y��~y���S�~�-2�Ӂ�qQs�D�L��g����/E�#��s�2}��D]��h�E
��)s�ޅ�ۢX�@�>0䞵|,��A�%h�..��To�
�7H~Y����:�2�Ƣ��eMQ/���k!��n�c���f��C�Vё%L��gv�x��b' �p��m����S 3���um��� l����a��x��1�H-��ξV4"dW����c�<�����%h�����z>P��p��n�ql�Lc}�\<��H~����Z��l0����K��(b�!Ry�q${��m;�j�&�%c�Uf*�ˏ�,�l�$���P*R~��oΠs��l?y��!���Q��HX"��sͫ��n~i@Y�S���@^��l*|$���Ɔ�+���x��B[L�R�y��?�Sm��_�N�S�[OT
���3+�@۸���7B����n@-	'�>|�i9v	�|�O�ڄlG<M��>�%5T�!�+(�j���Խ�u�r	�9�Yҝ�'��Qd�(Z����T�``	�/�Nʺ%}��߱�
����������Mc�e��	��6�������d|	����15�i�i[�Լ��˺�%:��g}:�D��'�z�7��cf;T��?-�i���$���C�7�\hp3�~σ�IW���x	��6Ɋ`������Nf�*�wk�Ez�bA�t�� [�#�c����2��YX�S4!R��9Cc_�B��7瘨��t��Q�
nG�=4�;R����S��gh����2�q!��NN��i���{�{�� &���N ���*9������A��ɵ-�E8�������U�-\��1,�mf�q�6�wR\9k�P��ڻ����}�TQ���y�)���0-qTb���ܳ�U�n�q�j���θ�MQ>[���5�����a��rH�� >�l�u�gR��C;؝����F�R�׹�0�A�r��O�B�
�580���CieW�.r"+ju;�H�뙚k������(���H�!���]�����n����gT�Q��\O}0;�@\��yZ��w��9q���7�6r�.2H���ў(��w��Eb�_Chf��\�f�56-V�����~� �i9�~z��h�"Ԑ��ϫ��	��������z�ȼ�����^�~�0�@{2�B0�9�T�?\(&Yi7	],,�������q���Km}FP<��`7n�q]nZY�K�[|*%��
ه�YL�]Ww�����Ɲ}*�Z�7�2&�F�U��J�o]�{�G=/�*:��ڤz|J{�-�]P%���Ze�O'�����T�#7�ٿ�Rn�z��(1�Tr��s�Z{�'h1�Q�s��X+8jn�hG�s�AP��1!\�i��	O���g��g��^;���8 �4�&��0�a��ϼ�o�lz׷�|��O��h�t;���ӣ�ʃӞ�p��+@-���7������%Wt��~�����5��6�s\�|��RZu�gAE~U�9���$��J{:��8�˪��No�/��(�@i�8��7-+��8��s��څ�C�����o�v�1��ӑ����3�/d�ʘ�D�kd,��m?���7c<H����{P���6r,���t���� ;z�,�r��YLBx��d�Ck��)J��IV8�b�qR�f�ez���Mɷȷ����N��a�����o�Z��!�"�%S��X���l3�>�?G�Q?^\L�ܒ���}6�s�3
�&���"bǒ}<d\AK$i�.{$�T{[�1�"X�#?(�-���EOK|x�W�V!X�X����g�9:�SAR�b�
��A��A�Ϻ%�D�;�t�,�����賋��g��<��5������5��&�1=���ӺVu�4s��sUiR��o�y�
�-�T,��(p�'�)4��SGF�W�H�Z� b���1@�����)�(R�}d�p��"x��E��]De��ʾ=�.G􁴏|@��Кw�]ٛ�a訥�c�:��D����lQ�]a���68l���h��+��ӫ!-�@�3�I�E���9k83W��)��)6 �Q�l�J�g��]��t�������m.N��GC�g����QB���^�:loYjo�n�`	�T˒�i
g�q�lƦ$��k^���ꞭＶn�m�Y*�l:C7#�E��ٿ6R���B������P��}<A�`�آHg*j��i��_\R�*�4�N~�#�H�E��">W�5�xJrE�F?�8�|���]f��v�O@��9�D�g;��]��y�w_���]�p3;r��{���^f�`��Rn���u6�*�SE�0����4./\������Cz�+�ڧ2�a��9��V�9��ؚB�}���O������U�֌�(��w=�S�/F���_�gM}ǅ�+?�001�k�n�{���uŪ��$��66ؕK������v�K"D�x�n�I�J��"��˴�U0�RbӅ���f-�N���������E�E��g��H�V�V]���^�3��ԧ��R����$G��⸎1jx:q߭����A=B�z�P~��4�[������Q����N'f�i 4[9Znذ�V��C��rw��#S�t���h49��{{��_�b����˻G���l�(�/���X.��������<�!�0�&��&�(�
^_�Y�|�(-|<!FW%�BD<3�:	��N�N�纛8\@�M����ўW��A���w���S�n�6?��W�Q�u�`�J7��� q5�z��F+,�R!��_=�"�hI���Q�7�����4G�e	���_�Մ��ꘖ�f�8-����P�nU�(pc�B7�d�v�����F+�1"Z�lcC!Ռ�Q�<+R�fO��+��i^1�c2t
J$�P�����w�X:��I����z��y"�~���KӴ	_y���o�w�6;�85�OF����g+�/�� Oo�A�0<c�К���ےɕuĮdsn�,���r��`��J-�ʿK���m�{�
������Qk�cF��o�i
@�Lh/nitr��NGa�����Y��xn����"����1B���6&}P�����J�F��~�B?��y!�Gf�����AWL�T
eе�ģ	|���҉�����?w�,/���%V���bu9��%S�U���?[��Q�b�=��RooMR��x�G�n�U���#]��Π�G����~&�ϐNܮ#�ŷ^�4�pI���cZ�A,�����g�ѕ2X�lPX�Y�`�Mx_<�6�P��(�w荠Vc��A@zC�o �G]�&��c���0K�5���|�����)6+����̀+j`H�ќ/���=p�)�W�1K���W����6�qE 'Nx�'=��\�[!cg���9W��/�6���Z�3^���{ϴ�v/��ͦZ����8Z���@�'�2�#3���YD�ɳ�a���۟�vlI"I�cz4E0u�����A�GҚ��E�X3��o0�WM�61��*E�F�����dOUy��8���[�객�Ւ�$���[��t������v	�qG4�-�RNP�-=-��H���|�؂y��U2i�Fw[U�rL�ۖ?�S#���9��t�A<�g����x�2�=�Q��M�=���N�aV^���M�ԣ�3X����]�B����2>-��������M�&j�|�08�ZfDH�i�o���\�"
aR����M���ܶhL��Bw%*|~�8O%��9�wD�{>1v�YLkIT��]N�bƤ�16;�
��=ë���y�K0 O_;���`��ґYZs���Ui��2��g-X'+"��߼��8Dv@�n��(x���7�*�aE�ө�cڨ"�#OuS�7�/�qaE�yŗ	�G<�!�a�O�0�mNXSp\��Y�ƣm� ա�l'l<���8�b�y4�b��p$
|�hd�8ʀZ�,F��T�"�p	�����PT0.�5�He5�m����ɤ�y8}B`@b��,�-? ��z��S�0%����}����?-�i�B܌x��x�`I7�&0��	��4JxC�kt�W[�bQ�],���6�Q�G)H��F���{ʞ��y��JD��R��+��r&����
�!�H� ɧ0�}�Stŋ�e��E���������k��2�]2��@w��C�IM
���Mt*S��K�L[�N�+#]���s?=��D����N��2� ���[��R^3r5A3f%a������X��g���f�NYs��B��,��_�^��muL������J�ǲJ`�H�V�c�i�Q�F/�'d�����ɋmv�]��R:���g�	���'D��xؐ!����9��%�LriK��S��4��\1�σ��8�w��{��k�q{�y�E�zQ���S����)KvJv%9���!(�	8����H�!��������#j3�� ���Fi͵�a�6�2�A�CT;�FF���ߢ�x���`X�����/���or-@1��#�a\���A���	ܗ��4���7�ˊ߁��n���A V�n�S��E��B��?N���:�1c��I=�/\��G3U�S�: ���'����+gA~<z$\�n�
���)��*�kL�3�4��ҏ���	u�ꐲ���FE᫕c�[$�����V"0��~��,��A^(2��/�'��Y'�vA@mʊ0��FsLT{O/2G2��,�'Xq���̝{��׊*j���(ǵ��Jmj� ��W>�(l8��֏}���yV���������_"���E����e8H�����
9�</���^*e�6n�a�0M�U�R�z����+&��Y��%���qpTşi��\,��_�Lh�E���SwH��F��*FY�sP��m0��I`�e�4�f�"\��?�?�R�FN
�6'5���/�$ A�2�a���	��g�d�w�z��l�f��[��j�^,~^(�J��HB�\��m����|R��]�ם���o�蓽dq&*2�X.5�ݗ�c,Z4����9��]�
`C��;]��@-��$�˩Fpd&A4?#ޞ�s6w��p��e�� �!Gg�34��3c^�}1�E�-b}5c�����/R�M�~�E�Fv��p��ɪ�'="�km�s)�AT?f�o�����}�?7�OD���J�H*1�%�p�=X�/�c�aZ���`�蜸�O�JWO�,�����:��	��~���k����C��_Mў�*+���*�D�R��Je�ݝ�[���E F7_���6N����CC�ĸ#Ǆ�f�
? 0����7�l�A�_�O\�u
O 'i�4wo��<g
X��i�<�T�_Ow���S�ѣd
m�(*C��R�QOM��m�G��KrS
�Vi ���xЋ�@�X	�xF���u\7���Y ���/"O��换�9�SZ��ou�lI�C�����%�αHz�	�x��=���S/]�B7�Lk(,���F�yܰ1��d��Y�I�8ol6��@��H�2t�����:��rucV�O�M�#��Q��i77�,(R�)7��D���D�	4�5�X�~�$��S�svE�f�f}���v���ݬRם�z�9h�*요:��r�B�@[�2��gCOkS�f���E����0I>'>$ʸ��}a��3M.���B5���/!�<������f_־e۰��%	R�
?ɥ�ΰ�wG�A�Q,Y�'�T�`������������2X�]�;�J�v�!q�T�~�bn�@�XlxVHYEB    a3ac    1230HN��kx]����7!�z���د(�z����3���S����P_��cQ�cE�Kc��S��K8��XR�UJRd|@wVU�=��6-[�x2??ےS��,`\��N�'D!9a�e��C� ;��Ak�u�U���E)xOkW�˒�׾�����I�
-���w�a�U�̢��V�^��?��<������IV;���@��!k8`:,)�f�	�����qf?�W['f���[�: ��+q����N�nE��o#2׌�mg5$���x	�g8;H�*ݱ��;�mb�%R"�~z\aX�<4��/ǜ|+���>�D��]r��Xo_ fv����n���e8�#*,�Ӂ9 ���"�T=�a%]3�
&�wB��D]{���^�Yd��BW0�a�S Е�KW1�fI2��\w7�Y�#J6��W��+̊=�O ��I�F��/�S�ʏW�o#�=˭��c�=-�`-Јf��К.�*�����T��������UH!t]@v�-U�@��Qp� �5�W]��(�x#ٱ{����:#/w��w�A ����)8,c*ӏer̀|��������=�?���ee�4H�t��~�f5�`����鑲��f�Fҷ/Y-�s��	���/�9�O��[�j�����AZ����ִ�}P��-��§9	����c�+�jV���EXY��ID��D5�{��y��Ј�
�(-fjd6NˬwT٦���7�(VG�b�5Бa��q����By��C�[U�J@���	P��Tѻ��{=Lw_$i:ݳӷ����Q}�wo���V��%�Ӌ-�m�Qf������pn�e��0�'0���"����h'i�V�"�)�@�-��6ŀ��1(Wnf�F�����@]���ͱ�?��0[`��DD|�|Z]�����q������u��m��:jr mw�%��ӂi.�)�/��>�/��z2m����F�[ V���N���K�9���"L=L���zZ�NA'��/�|��Li��%觤D+��R*�&�k���T��[l�~|�a���DcT�ߗ)�Z��QR�b��/V&���ܺn6��Hi4��ڏ�Ä�,���8�>���/���t��lJl0��@ηh���UB��2%{#�Od���_���t���V�s�/���~�<�0�Rw��U�w����{�qGB�b�W�Fqt��1.lhO^� ����JH��&l���n�3<�+�f�ߓ.?D�늕��T&������*ϛ+��&bF�>kG���g@�0����dd�V�B��C��s�psF�yh(��E�EJ2�o�ns�R����&��ç�<2�+����O�`�����U��'oi��ŋq�4�@<q����|���t�Lk�7�-�31}Xo���l��ވl�;@8��-Q������Y�� eX�H�-M1�����(����5��E���lGcE;�S�z<�A�Ř�9G_����an�mO󫩈z�x�s���#]$0��<�����A�z8�}#$�� �#��9�+�&��Fxo�����AiK�XWFj9)}�l��v���H�2��l�b6"�N2�7��X8��;�C.�
���
�Jt��ӆA������<�Q^gm�M��ü%ѐa�~����m�s��}^�wV�f��Ѩ�D2�uW���m����I5�N�u[D8x��Uv���1+�//]t�|�ыu���RRM�����V�f��Շ��z��HS�:t��W���OR5���1#"�\����bn�P
�na�ޏ�A��c�^���LL�_ɒ�ZL�K�m�W���7���lo���$s�����V�n�Er��g@�Q��6���.6AXnn�O�d��Q��W�=n��0���Ik�ĥ���B4։�Z9�0���)l��*C1��7��N Ѥ�	�ˍ]�5�EL Un�B �zmʫe��Gͣ��Hj1ݚ����
���>�O��>�V�+n&V����Թ�R@A��@�����4˒�������bB��;!�x�A�v�ZnQO
�`�}:T`V��0��t�5-���� e>Fl!�����vv �ҕ2�º\���Ƨ^r[~��(H�D���0LOu�j�,�w��#u�bc�E=�=�`� p�Z�%���?A���S�u<2QI�'�xo�O�?�s����Q�Ơ�q�7�ee�CX��z�VP qm[g���i�0D^*��v�O�X-<��9p��81�Hq����)�I�wU��_y��y 6l�*����~��?�,�S���-k���WP �ds�.p��U=Ц0�@�S`�G��Ze׆���YPĬ����r�����}�����BQ8�F��P�zD�g�������d]� �˼O�1
h�rL�u�8[�g��;��W5�(�\���_����Hs�*�����=O��3��)���}����R�钌���m�֒T���䅣Xe�@���ӗ$<��ISQ;[�w%�<uakDU�[�ԢG���f�OޮQzdC����U�0��h;����E)(�p��3٤gzS�p
�͙s��F8��u&^���K����ןGp�C1:���0�BX�^��������y��v.g�*�b�P���|�v��?�'���J&@�Q��e!i3����{p�h�O�� ��eἷ��V8A~���H�3d�g��%���X�8��P�����?�ø�����H绦.�03	ͫ�A*��k��`qo��	=�#�Rū`�Q����m#�LI���7��G���T�`�u9,��b8c\���$u����^��\Z(u�������c��4�����/K+��7hU�MALPzH>��U�7޾��9�Q��՚���;�Sd�����ˠ�O�$e�x�d��K��.\��PP�ц�����	��k���|�G'֒Rx�iV�+��b�Д0��`�:p��w�L���js (��+���Or�hc�\�}Bs��D��w:Q˙�T�����n�w��?�1�nf��P/9��J&V�����5������.�3'x�y���>��̮�p�DQ�@ù�i1��8��*LٶVڰ��!H�a/��)�T��31�tU��/�LJq�A�����#@q��TE+�Ԉg����E �W��_�����ш�*l��Xl�E�ہ=b�[�&�Z��;�s(����2�-Cm���	�t����ZDe��.�Y�C.��&إ�C��$I_�e
Fn���WS���0����O6W܇AqL��(D�0���^�Ef��ke.��l�-MJ����v5�� 
0W�P�B��lp-�$��XT��I"V(� ��;Z���e������8�A�	D�������$%�x�c�;uq���	(����)kx�>����9Ms�|=�aP��H	��^ [�|�sneq�::�l�@�d]�2�jx&ՊGQ�\���1�x���4r�H� o��"K�B���b���L'l�����ۧ���k@p	�js��%�8��HR�3���u�W��[�ԓ�Wכשz~ALҖ��`ra���'0���x��6���JP)D��ȋ�>D~N���>Ě1_�	c��Vƃ���c�3��Nhn�Z1�a��"������kt�='�/ ����uM�;9�'Z�=�z��L��(]tl�8Vt˰�v���8i����L�������W�kl�oRM�c
q;?c����8��.��w�o5H^*��(9AS��w�ی��I��ݞT�vcb���0m&*dZ�zg{uO���t-��H�v*����nT�/�R�ɱgЄ��1�#�[;�ҙ���c�0V:��3�3�&Ƙ���u4�`�m�O �#�-�cR�N�+��OT�X-$Uĝ�|K�.\mp������[c;�p�g�&z9Y.ɦ?a�lG!=ӟVF� ��q�.Z�Z'Lp'�s{�a&�D`��x���ZIy%�^�rb4�/��+)��<�"-Ե(��J�d�wV�ti��{����g�h/��rG�X{�y���i������K��y���2&�J*�Y�ua]3Cgx��R*l�%@Gù�w��Yى�,��2w^S��v1��Vi20��/%�`�v-Px��f$~Ik���u�9�a	N=!<����!����"��K�k��\m>��B~��!�1Nc�rp8��if�;^�~�62��� ������j�MHEz���x�/�1��V�����nwկ�w��>b�v����C2a�'ak�$l�>��eә7���V.���6j��7%V��$/�|+�@ 9�ac�A��T���}�z����+��n����i��8����;Ŗ� ʻ�}�^	���Yv���~^���m�P@0˲��G9�� �.w�����'\��K6�oT�S\�T�<cq�9G媹2����#Z�S��w��-��=Q�!w_�j|���!v��G��10#��������o��ߜܰ�_< WH?KJ���>���~*YH��@շ����4�;� [Pl�㽌�+>��<��`ZaVNHg�p���J�^�1\{R��w�ԙ�D�Vf�	�ʉ�l����ٶ�ä�� 5 A�6�)��