XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i���j���9������ �����퀮�6m/�
Æ��>�h�I���Io���\�������i�cê�k�_ݚ~�凟���چ�0]猼��>93�^��R�F+�^���&0�y��a�Qz�/`�S���.f��W�2W�S���{�N�P��Ծ:H6oA(�^F���M�1�s�&K`ut��ǌ�נ�i�+�t���7Q�.��,'=:S`i�M��9��abv�� GϜ��eߚt5�yl$0���7�"k�bUz-q�zz�g�	��rP��wf�2��;9�ih�N�ܠ�[�?��ƚ�P���ǂ,�`���s�:�uؔ+��L���t� Fغ+�:-�xw��F4
#��)b��Z3�d���$��w_�<L�~~��\���;H�����t��l8������ڶ �3ʕ!i���esK\���<����$�U�1��m]C�d�|���-HZTu�6;~E=�3��ɍ�p�.����<��Y@5�Ҽ����cc4��̀�����y�*�򦩍�l�	ntF��)���5���/B�����5��b�c�kO��A?���r�1��>+�����j�OE�r���M�y�(�������Go���?��S��N��S�-}WTh�v:7���K 09cX}��{��,��`3���,(]	i:Ў��u���0�������M!��u`CJ	�� �(6��<9Pp�8�dm����ik�]����_��@�)����k͵#��t�K��[���>XlxVHYEB    c3e8    1d20�U7���қ�ʎ�p��³=�{�������[�}E�Fx�p�'��{����-��F�u�~|���� �Vƭ��=���$��6����	��9	nr*�۠1���%½p�C�L����Ϋ�c ��/]��|T��u����"e��B����H�nO
#�tH���n(�pNF=~��b@��Tv�o�XӶ��!Ç'��p� ��4#y��Y��fI]�����ӵ6��ڴ��1Y�s<gC���m�`�u�Ґ#�K҇;��X;7EsF\���'�5��Tr/_�x���5[�RT/�&<�Ci��������,��*���-~�"Y��U����j�z��Z�}�go�C7��O+P�Aܬ��R�n.�Ȋ�}n�x�iM!٦���Gd9�����%?��]<W�B �TӰ�}c�UT}
_gr�6<�hY~��\L�~u���/�[��|G��A�������P3HIl�:<+%ѝ����霵3rٜR��%��(�O����|@�q-�G
�v�z�.1I]4V����߰�وɍ#�=:�_�g���y��F�Cy���Z����2���7�و�0k�&V�хd/1�6��b��}x|�p���m �Ɉ�ֽٍ���w"�D� e��רּ�f���'\_��Q�Bcf�5���L��ڠx=�X�.@S'X��J��`_|�.�U�rvð����6`j��`@@*n����xk��U+ 8z��N�F�,@'�ꦀ��Մ�j���o��m2=��^����2�	�ι�p �JvH��42��%�F	`���&4ɶ�&�8z�z�X��nab[L�,�g�|{�ͅ�N��SNHxg#ox"6����p�>�U� ���4+�yRI�����ʎ>	|�;/4�{�w8|`a3�\�6�����ZH�2�e|�{V�Ti;��������<���<*$څ_��`������g�7��(��]ׄ(��![�y��ѽ������f��*��q���4�$w�]���UR�9��>�����Ti�.6�}���d�_�	r��|]�#hј15��a����x���`%�2���Tp}g��������HZ<�qU�C���-��hn�"1��G��vL��xTzX��:�����m�̘��$�sx��.��Y>ADs��χ5H;V��rJ�6O��r�D���`c��>�W6	k�ӈ:��l+F�( O���5���U���gl�w�}�U�������K�H֯��R��ZIox�rJH�~� �E���jb��v���%�1�J0qk~��C��m&����خ�7��~���wuj�X��C)m`�K/�"��Z`��N'�eu�g.4�Go�|f,p�f�!��fZ��<�8�K���C��2#2X�g-G���t|�:�Os-�?�c�Y%�������3S�~#���I���A,�f��iC��m�2��~���@�>���~��-
�M�l�[��G��rjq+����YѢ���9�����j��(^���;�7������ADl3���δ�"S>���ba����~�y]�e�h������/(�2�r�c�䣺��십��Zc!��YV&(/pp�"Q�;��9��gHӮ��"�5���0f�2�Z��ѭ���d�{?˛��;Mnm��~r��mM�BS��0����
nڻS�`TW�P`7��x�i�
�a#<!#d�I�}u%�4� T���"��`��H�Z����}}݇(�E�kXo��E�
Շ���2�4SZ(��dB6FƯˡ!p��C��݁,l�h.+�� B[#��n>�س%@W�d'7;��������]�A�׌t��Z$�xM����<�w�-��a�L�cz�K����JkN�J2����64;�jP���� �Hm��^�]e*�Qv�KaK�F���'j|N!���cXlb���G;�Sî([X���>MG�E��Vĸ.O�*��ǔ�w�t��I��sB�WRtV ��i�_g�&g�
��teI��6b�(�a�݄#.��=P53��	��2F��y�Qw���mO�}��,8	�����:I����CS�oGH8>o"�D��%r&?a��<'\�b�)ð�r�W)�]X<ysF���b�K}�\	^�}�k�S-_$LJ~�|ڢ2-�u��',���p.�}B�_�_�s��Ж���%�-�/��\�88����&���o&��BRp�Fq\
��=���-."b����Y��
=�3�-�CBm(�#��_��a���[�|��;3�W�B;�d�5@]�+�G����-�@�1�"�S�8uvW�KG�������'�:����ƝrMyQ�Z���bi�{L�jOpR滟wO�DB�΃�b�Ө��W2�w��x4�f�}�
�?�D��gw�~�$Z�>
.v��&� ���,��?�艤���Vq�]V{D�s��O�t!��f%Z�E�y�½8�@%5.�N�^aɖ`-@�9!jG�<)��0A$w�J�°�я�D<@�L��FP�yc�%��Iq�)�s>#�Pz�=��E_���v+�7��*������`�W��*/A�������c�C�N��4�z�Şak�`�E���	B���t�Y3j$nH����œ���ç���_�IN����^)잀�U��Y��DL��^K��b�W~U�1����0�s(6˭�c���E�iv��` ���kE=�j:I�A5�Sx�!����ɝ��,u֥�Ny.y��eJN���n���'��t�)���lz/�d�o�h�Ne�{m���� ztCT ��^�����ԕ����Z�n8�|�&��I���V$���\*��q^($(�釣�ȥ���U�--m��\�X��o�O)�Z2e�7�A�T	�mMbu6���C�@G�ꄤ�"�?�9[|,�G��$s�,'V���e�f�u=!AG��nf�V��Y��)@"sՒ� ��㏙���{��x>C��c��e�/��ԑ?^�PVIk(�py���>�� �N��'����P�;�&"��K�]�dZl�a�E�u3��������ؗ N��>8GX3�y�Ϗ,��P��j��4=��Nx�q;����*N;A����g]�����ӳJ�#�8�jP\.�����u<�w�x�5\"`.�D�у%�<�"�Q�� ѣ:"�덒Ʃa�]��R(�_��h�y�>r+�l�S�ӂRCjqb ���~�"t)s��*���E��\Þ��b��&Ȗ#�����c2�Ou�Okƕ�&xs��/�~��t�d���yۺs�b��v���X���|ˤ�s"g��f�:U��)���I�����U �{M[X��B�	͢m(Rc�/�q��:D�?� ��2�Y 5�g�Ò�uo� f�]��fb���<u��=�Bv�T���u^A/��[E���������x�;瑳AV�.�N��U�>Hj�ӽ�T��:�(��`彔��p�����xS|W�$с�t�-<i��n9(ch��U	78+}~�qn|��US�-J���XٺF{�Lt+BA�?o��e�zj�d��u$�m�pmb\�Țf-�OK-;�п�u���o0#�yz@F>g�2�vd����s��NGv�
�2|�T� tK�̱z?.����b��'�4�Z���l!�7���,��*�.��]��_)���i�9y-��6Sٱ����9�����5e�͵Y9m�*�
_�3�l0�eT���TVE�A�����LgH��\���%�;͌f�Z���^&�X���1�P�sw����I2�6��Y=k�>Q��������6�/FaX�-kIz'g�@���O�ǀ����o��+3v���n։!7��"�]+"�s%�O��+��4u����%V��l�)������A,َ����);�}d^d�2���-y
k�9�P����M5�L��6�& ��	<�Z�wtޑ��/����� a��Q�U����Y[�,���A�K�VE����H0�׮ &6�mJ����uL�';jג��uf)2q8�ɃDASYǄ�ej��u�b}qZ˘� �&Y׎�c��D�,3A_O�_�*���a_*'))�����D����3�����|8�p�׫Y����E�H��N��jb$23-ւ�d�����F��
RS��i��K�-�}�2�L0�ai���4�x[C�q%[��Z����9�&�%_!T�_�.�U�Cġ؏Q���t�Ϲf���<'p���{���
])<O�ѻ�_`�<2Ҷm�}fw��N�Ū��Aqimj}���#�k��e���UdD+��N�!@�9�D����Q�tJ�G��$+	7	������j��{&о���C�֕x�Nf��yYrF���	s��&����!��� |� ����3��N�	�}�2�!#Eo�4C��sE�ø�x�0��x�d�ܯ�Ke�EgF�����e�>Q��,���W��,�k��xK�j�� ���p��/(媒��5x]l���VW��{�|����z��t?�OSr�a�ʛ���KXæ���x �u�[�M���LA�U��%���J\tx���3.�H��}���{�(��rt��������{�_\n +���*˻q/��P�l�HVJ�����S�"hNvd����k���ݘ&��bJ��ADu=�d���%��O��x9��Шn~��t���6�x�3�9yb��11[�j|���en��������=��j��D8��A�Å�[7�Q,_�o~�.,��z�����&8{��.K���+�޷�hԵ�I�,z�3��e!���<D˾���xn\�bp�z"׼:����i� zP�����$�{���֔�����߁�ѿ��7̴M�,9qU=;�@���������A��,foT�q4?�J2�^U��08Le��[m��9�$��b:��7����vIFU\�RiW �a����P6�F���-�|�\&q�Y���k�6S3�|f&Ψ$�6ն��5�<{����w�]�ﺥl�4���������ͨ���b�"�r�.�}wѢ �re� �pf�����O����c�)�򽸺e}]h��,�gm(Ϣ�hZ�p3e��s a���J��$a�+2���7�ˍ9���M���:'�u��}���lC�%�g�	���({���:�k����(���'�0��6D���7��%�kCI���B�P�w&x���F@���ɳ%�i9��`����bp.�X�7��)	JVa*���JZ�92s�E�y�7'r���v�8���4O����l]I���DS���2V��#i�&/�4=�/o:Z�BfЗ��^�&�l��T=��R1&��2��\��U��/�����#�O��{ƶ�"��,p��+�\�>��F�N'�$D�~���[fʂئ$������f����X���Ί�����(��i ���L�"u^�[Z�J%0�]�G�{b-��13��p�:��;��^?\�����䝶E�����{��g0�X]�4NCjL�ie*L���`?�a!�>�[9��/m��^�|��=�B��.�5ʪ��6칋r,5B���.3lS�/�X�W2+��-�zS�̤P�_���~��+�f���ւ�w";Oe'B�	����0���P��f@�hz�1��+u�.�$�e�n�81&ײLC��QV�2679�C���2#�m��G!{���ʞ�_J�!U��TSމ2f r�9|`�J��D1li�,^ݡ1s����/t�W���t�o�I|�-��0(a������#.� U�Y�N/���8��Hi���Ȣ<H�nb)�2p��"��QJ����<b�y�S����!�ՆKX�s/}v	3]�D��S�Lnw�ៗ�!�ATFaXԼ���$�Q��d
�M��v���W@$X�Uui�~x����z� w�EP�}R!c9���C��o
�>��耵+���BϪ��HL������o�O0����Ӿ[k����ga�P�-�s��b��a�]��n{]�e	�F�ùuB94���+pF�@� b^��f M�Kc��7�#W�tT��vԄl�Z���d��q�]
�c��?��R�~(w(� F��;t�:ό�x@ڪ�K��U��dOtݞ23�Fи1Y��s�k9�I�mk�v\s�Mc���˵9� ��:��ynL�9�tص�	P~g���{��0�C륽(���h3y
�9�[�{���YT�T��RR)�C>�wצ�`G&��&!j�d$
o���k1G�̰Q?'=���f�!Z4�_^���z���z�*8��"��}�EPO�SR[fH��y{�DpO������t�������̱/�x?/��s�����OΥ�V`�5�Dv���;�Y��P��5��tM����~���_{�6��]��V��5z2	�>t�x����h�t>eq菴�c^�w��x���� FU�ط~ �ҷ�D���M�	�t������ OE��#�dW�;]b�X�J:���#�5��wN�J%<�	;�5��<03��U�Re�#��>�9�j��RuJn��y*�;�Q�����t�FFw���)�*���b�?Q0z�;I��� %ͅ6u��0(�����*I*FW=Jaa��	̦�V�2����y��s7���Xs�����ٌl^�in�g9 �0����nj�D���j7�]s�d �TT�{��?�5}�d�!v���P���V�DP_��/��5e�L�6�$��7��g���'�(	��c���P�A�[Fl?S��?GW%��˫FW�0��WC�]����I{�WoHx����i��'�+�8��3��A��,�{��0��1q�u������E/\���� �0�ʜ�R�#>�iL �^Wec�#��ޤ�o��:���#��j������'�E-�\��u�]��r�^�a#g��A)�R�=ZQ��H5�
�5p_����b!���VM�����t��iC=�N�sڀŭ��R��ԻV-��l��h"*��n��Yk0�aO��#A��_�#�޳�uN�}����XylJ�
0~��-&�$�Y��~�+`~�D��S�.r#ڵ���H�V��J��	
�,�Y�J���}�9�B֒
:��y�H�(d� �����pc#�0�*�4-6sJ6�T�Y����L��)���'yϲ���n�������ٕ*4���<���}��5�v'm�J��� 9�X�諢;q�ie���VPo��t����f4u�Jy	[�^G氰T#�ޙ��*�h���Q�$(������TFy9r�V��kƀ�ڵ8%JrX��1L�Y���x�g�����|��,���o��3&�5*�GL��S���B�����xT�H�0��M�O`]�uX�������XS'���!_�g�