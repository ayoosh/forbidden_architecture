XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x��A��h�W}z�9,]��UV���|��R�pi�.���9\^,#罽�� �J���,�h��q�_��"ӎR1�����J ��^�?'��5��{�l����-%��.�ڮ|��M�֛�H�W�}���`�W�!��1������v���=ҵS�H�����QK���(��9Q�)'L� �����쥊���w���0�_ƏZS��c�Y�4�kt��:�ar���%%CW��2��,@��7�~�xCp-�r-FFGDK�$��p�d��pYe�H�Y Nǘ8�;&k���WִS�､�N ����G�e}a���77 	 ����$�ǭv6�l ��%J�G��ᙠ^���u�vO�6��`4ʕ��".$W>|��A;q�.��G`�c���b���� �EQ��S���wȰq��`[r|؈Msp�̮�_d>X3[�J��E��}J�I���'rr�*�ns��R���ￒ��4�&	��6��[*'���s���T]�/����ŭab;У䗰Q�ʘ�R�r�G5�6���8�!��������aM�:�8�k��������"����
�#/�Ϸ+�-g���	1h�P7{m�W����Ћ=}?h2�� c�J���]G.|<;-v��u|�P)Ӡ�8� Aܽ��QVB���]���q�rp�����#|IAv� i�b�W�
U1���M�nn��6"���7{���rX[�C=F�h��M�k�އ;�ڨx�L�|c��p�❌�0��z�XlxVHYEB    c3fd    1d30K��OU��Xj��`v�m��%F�ќ��k����	»�s��]531 ���m�.s�s#��c4g����r^�'K#�Doy�μɐ�X�b;Y	��H�~�O~	fG�����ӯ��?旼 ���y�0=���E�%��pE�&X@℥��O��B�}�O�(��Ǹ�y�b��m�Ѩ�ԙh���c����� ��k��G���R�"ʡ��Δ�����&��J578J�fg��b��p��a�|F�5���#aYϾ7���γ������ �ԝw/bT���lJ��qN�.@M-�G��d�~$�*�}5�t'@�B�g��+s��KS��QG�#{4��˔l��ѡ�eyB��9�&��^e��C@�Xd����s��86:cw�P��)$�N�U�bz|ӗ����k��i�to�1�j�{��'Ե&s�q�R�X�ǣ��0{���T���B'f�ohWT�T�ЌD�w��(�/E�HFD�2t`_���N��f|��`�L�R�
툦8cG�蒁cפ)ލr���5 �)��@Z�x��;�(Ka%˖[��p�RX�n�D�q+{}�6�0��
���Ǎ�ݙq�^�� 7i^�}bXY":���Yɧ
>��7�p�6Ý�ĳd�E��J��.D+���sE��6u�{ �Sf�2zw�Z�W!��OY�;��1S��h��mJ��V��/�I	W.����JF���$x�8�.��z_Jy�CRa߱:� 6�3���/JW��shQ�b^W��6Q\�wu7���w%�o��h���ۦٸ�ll�{��E�"�-�̳F��pUH��ʐ�7���Z�Vj���5��1g�@p���:(�4<Zv2bH�y[��d�Ě�u��FJ,�da�h�BS��㩗�}�Yɒ� ��~�o '�PN���	O[]9h���>�d�( �:K��"��R���p�tH�����w֟+��|daWÙ��.��)D5�oк���4m�M��]�w�"Ť"{��m��>���t�B:��=���IRx5��d����?�}{��a6ۈ�3躺����|��2A!>:���C�^��-:��5�3$�Z�����2 B�M#���JT�[����Z�p�fI,�[�t���~' ��{�n��@�i��3S�.����AI\ϳ�1ۏ�!��c�/s5a?��),>���+z��M�_��<�h���
���;�d5�s�!_Vca�Ȩ
���T��Xx�������+w�}��|JJr�ko*f�
�w�[��p҆j��̼;���ѡ��º�S�3��)���N�Ͻ��ǉu�p}\��YP����U3��̟�
K�(��kA"�c�z�Gu���Mֳ�g+G\)��:;j{ğX�.9�-5�'o8{�<;��E OC�\ ����ہ���O��<V�e�nw����?�wI���ղ<5�k�C� �dC�+c/��?�~�@�#�E�Pn��%�X�Q^�ԋ��0�
w7Lq}�����j��/�;!h^���a�V���<F
ĉ���Nk��A��������&�|2�u+�1J��Ԥ91t�]�w��0dT�9{)n�)wH~�ٴ�tIB5�����?y짂�3�Lfˮ9"��mX�0l�{.��@jJ�bB�riD��Xuƾ��"Hs����M�J�ԇ�Q�� �Z�k�i�j��	��̑��1�u��^��٫ȫ9���ք�p���3�x��B�&Ŀc@����H@U����Ţ4&.V�ĩUG%i�^G ќc��1�6��ͻp��o�����o���-5*�b}���=���~努E�Yh����Y=E���n$:����ݩ�yE�;���׮���KV���ߵ�J"1(-#oETT��t#�������U!�.Г{!,����d�<H{)�K=������b�IvA<ҼG�)���z��������z���������N8�B�`!�o�l�&t��I��U}(\��&�q��t�B�n�u"D�v�F�9G�\�D�2i�|Vg}څ�nٚ��?A	��an�̗ұ�����G�(�7!&ڳ+�2T�+`أ3�P]a)"��k����_��R<Y�|ՓGi��n�`��B5i�R�R��P,��X��b8�s�����ֽqVs�F/,
��a�Z˯{ճ���oh9!<B�o7������l}�$^�掣�w�� @�r���[lb� �à��6D�;�2�h"$����vF�UP�_��r_6��p-F�x�)�:�,\�wG��i��]��I�P`���z`G����^�O�Ϫ�y��^��`�����7w펕0nz��XB��eF�}�F��cK��B��e8�K^>x&����JdؾJ=�Ył����9:a��^\��7���4s�1�#ۚUh1�ڋ��q]�v�!�C��c�e��I��A��Dr�]!�7��������jcF� M6E:+�_��`��Q��>��Ƿ,�`��G��
>��&�䅇uG�, �r�3��������+ T14�R�ǵFi4a���C��e|�7%�����8*���̷%�6u/�m��h��]�L��8��R�{]F9�tsB?�(�����_:��]K��yT&�THN���M��4<9bん����U��+��/j�ܜp��a�z���롙�"��|*��B�7�n�u� �oֺ���1g�. �UA�2�mS _�ׯ!����!��G�0A�2	M��3�{ yPKM�ܫYjĊ|g��I��.ԦL�D��sꍚ�0����D���М#��9�����I},C��*gB��]��?��5{��V�R�e�����|�>�����@מfy����[�M �lX�~B�������74��h26�hn^�Q��̈́#i�J�w�,a��ݕ����*I�(G�7l�@�����F����]�Fjc�C �a:�xڗ����J���P>�t�$��T?�\C����f�/��W}mEJ�?w�����͑+�|�$���ܧGS��;�x�[��Nx�Ȫ2ؠ�`4����!�3D02���ț=�?����W���=�^i?&����)��-r2;hUA�l ޸m$�����M� �W}��O6���Z�9jN��zD��*��?��ǩ�u/�M]�:)�;�� �Pq��Kv�Q��VRj�`��j�kF��*�"n{\��]�{�X��9#s�-��/2�V��f�ve�@�|�bc_|`IvF�-5���a���"Y���s���re�+F����>��+��;xx}��[�fȒ�ۇ�F�r�;J^��s�[�:M�2G�H��}��CX�?}w�	/���t�[�j�]�,e�vR��+�C����x0����t�u���_�T�
c~G/����P�	�y5�oB����Є��� DK
�n0s��mc.��v�Xĕ^�P���g�����Q&����*�W+v����

j|JaX�°��?���*���Nxm��f����v6�,�}���k����*�;�d9��oR������ ��Q�1����(g����ӻ皴?��s�Z8 "�޶7�G���8��k��t���՗�|H�t���5A�D��
n�1�Q�5�P- Vh�	����6�B��sE��DU�	�]Ո�MT��c��u���9���C���8�#,uK=C
=iQ��ͷ�R���F�i�%,$�n�$����U���w�����X|�p��iH��,v����6�h/�!�D��#\ }/�Ez�:�"8����Ĺ��;���e�xAorg�>"Ԫhf�����؛�)�
���~��Us�]+O�4\�����%�8nv^x���gԼ���X�'��Ӥ�n�T8ˉ��K�� �u;�5_P�야�7���#1�	�;I]}yz"R� �彠4���ba��\���Y������X4��7��"��y���P�ZD�°d�r`�Ӽ縢>��>�MRr�*��3����)NN9Zz�wKb�o���Ѝ�	��n���m�G iU�SdV:��;n��o��Y�W���AX t]}ky��$�m
���Ц�ֶA�0J���~�u"�Oo���Q��8"�i�Η:��!�hp}�����ޠe��ؓ����<��m-L���4~���!�=��jsƄ,Pْu !ṏ��Сa�r�]��#;Q ]K\�9��&�1^]��cL|�����{���������];����ޓ����e�| �)RP"�ӴLZrU��,����E�V̀t$L���L�&�^��(�X�m�,SL��Bv u{[�u��0��#LM���GՉ��X
��I����l���W�RC��$_��D,c���x$<li��G�Z�
l҈�8�d��~��������[eEQ�<!3r Q���"���xL�fTf<�õ;Z��儀!o�5��<���Z��m'u�~G��k8��l����N��>֍��O�!�F π��ha�4��|6X�W��h��,�s��5@��t1��1F�	�2�F!��!k��E�穆M��l����9JƄ���]�}sX�T��5�����}s��h����]�a�_�qy�5TT6�1x�3��$���}�i�#�Fn�t�y�
{��Wʪ�å�k�x0�5�E��vRT6@B �z%���5����aA޵�����s�.���)"AĪ/��W�*1ݞX�����ʐ>Jd��$�?� LS?�&Dt*��4:r�Q��t	\���w�\֍��ȑ �WĤ����}&�������?�!��Ⱦ��>:���뛾��:7����rxz������>���J���	.H*-�����h� MgQnM�^��BO�މ��km��9�� #��޶/�lU��P�(.����$��N�=�-��C�i6ygir��ķ��܈�z'e6��5��a�`���P&LQŷ�Y�~���&2hy@"���YE��&R�3�_ ��w���������8x�B9����6����Q��V�|���w5����f��
8m�s���d��"5"P�����"�Þ�l��<���^�GV�QZ���0 ؁x[:�����0i�˰za�k�� ���\��\KDLm}a�y���A��7�v�����������t��0�4�`t]aO�mz�O�,Wi�� ��S}�,U8n4=��`\8�'3�]:P{�<�+%��4�[B\e%��j�1�oJ,n�^��j:�zמi�C�ܥ.f�d��-v����<70XH����F̵m�6���e�{��s�J���;t~�N�^�&x9�h2#�����{(X�yR�L��zw��T�e>+���=�ѧ��6��n3^JX�8�\�YM�(�T��H�t�ݗmE\$oy�e&�^�7R�v\ZLXq3�t��
�h��6*t�/)`űXA����K��%�P�
�T���ڂ�u�a��=��9��Ѵ�̲�s��ٷ����O�h=�]�h;b��̕�bV��D>�	&���T�=4w;c����Sz�p�������k�1:��+4����~�ymH��e�{�U����.�];߫���[�����.fj��u@z��5y�(�B�+�����)�u6��̉&/�F�h��i�_a��^{d����g��d2#���˫��qo���a}"z�|�)vt�o��j��8���Am-Le���EèH3#���v��bK~�SH�+^�K}'�3��rח[>/-���H�
ގ?ZA],)�Ǉ��Т�l��(�u/1���j?�M�ڂ��AAI�Q朩t���s�1������@���	Y6�%���>�ህ�fc�ˆ�?<�����4gʙᘷ/xɎ�M�Īh�on��:F�g2�0�Sm�-y���EPL:��R�0�t/����E@����)8Jn�/Xu�����������<S|�Wh1I����J�����yS��'o���qn#q^��� ����Y�p��j�o+��d�
_�iM�;��2�c�g�ȃ�'�$������ʛ�I2��`L(����!(yG͊<l���<D8�nfq��Y����4#P�6�����V�a�}��ۭ%O�Ȁ͉Ct����R��F��¶�s�K�}���8�����)���.�J���7Bef�NnR@ �]�MB��m�?jK T��6�@&��&VGVi�׆�И!�[��[����@�V̕$�ND�u�K�9�'�4< @u\]�GN |��|ϙ4dUb��W��XP�w�/����dY�<�d��p^���滫�C 2@`�`/m�2�ES�i!��kм�!���~E�����dY+b��D0O�������r}�it���f��c�Ȓ�1a�y+�ߺtw�'Q�#�
��l��,�1��2������ ��]� ��eژ��W����1���z�5�9&b�wtW�(�,���K�ֶ�4	��0�le��/�������S�����уЅm�"!�\t��n��^��u����,m%�^VU�:)Cx�@��W�O��F�R��$"�����p�Vإ7+ۦN���~�n{�����?^v���Ef�B+<��>E㡾#��č33�
f��m�n����ա��~3hP�9S	M��1�3X}D�Q�D=X	zg�nq6����a�&jc���m"��n�yI��Хr@��́�2ʟF��	�0 ��உ����E)��&֍��),���(���^��NvO�;�5�,J7Ӎ"<���gz0�0v̨
8�%������ót�.���}1�=�U��=�n';	��ק��Gs�{C��|l��9c�@Ю�ʞ�A��>ռ���fwn�m���w����'�sѹ�Sj�}��Ȇ�e9e	�_~��ǉ���V��o�?�D�Y�V��B����~���^xge��c�X#Ӎ�zC�����G1�3L�rAe&g��ރ��ϵ+�gȜ�W���$ :�A_Cx�s�dz�qh��U����K^���!睰���"|�p� �Yd\T�p�2>)���WB�/�Y�r��[
�ℊ�����4�;N��"����b�9)Lуq>�~ҏ�����Q*�]���;*�n�s/&�$����#��M�~�������cɛ)�^\�zb�[�VU5֭��ѽu<c�}���}2{y�G|�88E���ᇞ�0vǛ��;��~؈}P�^W0�:��^ ޸����Ǣ��VN�(��EO܏�r(���ԩp�+<����aB�3Tk�)d �	"dq^d��6*�3��֡�,�J�{g��@TI'*F�}�����4OS'9^X�ŉ�