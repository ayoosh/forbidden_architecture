XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��lVȬ����A�#��T4���pC�t���R�m�(t��DO�YY6��R�Ӈ��;�9��
+ȵ�<�MõI �;[�T&c��9 Ҁ��;�`���@�ì����Rg��6b(�[H?X[aǃ�s�����w#�q�c�z��*ţ�E�&z�]�a��Ϛ��v��r	���D=�s���M$W�>�9��z�85[@@� .@I�B$֕z���!
J]�R!�ܣ��2;��hA*mGϖs5�������^F��9�"�5����i8k�X�C���_W�� �#��.���*�լg~�Y�8��%'�VM#�d/����o�27?`�4�*��g�'�]<rP��!4h39��.}���%>G@��]���C#@E$LЍ��iG��
aG��u:��&u!��Ý��Ķ�A��g��A���2B?��dU%@lG��C^]O]�_j�w,G�͟(��]UK�杅�9��\��<�X��B��j��
�]����9&�E�kc�L���~�l��R��`�Թ�N��3^�>mҧb4��*M��&���������	�JGb�G��5ݻ���"i'�y�r�m�&�[�G�R�b.,�am���C���7�a�������Ŵ7�p<0�)\F.]PNv�:����k�9���	tX+��ӈ�S"����aL�j]���%b
ur�T�VA�\.�Ea/�+��0���\)�Q�33VE6�'eh�+{���tr>o-¡4*�6�'��6a,�����>���<�{�;�XlxVHYEB    fa00    1ca0ܴ2����ym¸U��NOo&V'1�����x��#�?S�~A��>�%5Ý�t���S��Jmh�o�Em��s9P�pT�=}l!��	�2����S��K�`��#G��oP�^EU�bM�F�:s���٢z��z��N ��û�
I��*b2<��~��.K�e3E��]G�#��r2�f��m'xAOb5�M�yK��	�9�~U*Ǯ@5�r]]���:�f�wC��3�HƸɵ�b6�6��
d�>�Ы��n��m.�P�ث�,�ʶu�@�>S��_�8h'W�Z.��L�&̫2U(o��b�T��ue�z��>�K�%��^ɿ+E'R0)���4�T��{�Ԑ8��S��E�Y�L�'^�����D|>������D@]$k����t_ʙ�ܪԚ:7�6q��>O �U�x2��QB=��.�bC
[1�l��ǍV2%\-��7cS�����ɖT��Q�V����2/�g4��b����HL،�V����	�kc���B`겜�q���c${�-�5)U�B���3���>��}==��@Re���!=~α�6<��Ed�����|[#w��L�=��!	X�ʺkQ�^$Ap5����q�̄31O���h�����C������
�@\a��I�3Ӹ�Li�pL�	?3�f����r}Gp��I;��V�\�����V������-b�py
0����f�f��cF']=����̾�=�ñt�A2;}�"��e��UCT|�T��ႝƃAIe��K	���a���Q��v8~���v������WH�-.����������{׾ro�By��hY��+(mlɲ!��2C���<��>@z\�0D�j�7.�ʁESI3\#+�f@����*�ݎ	�d"�'�u*�.(p����&X|�r�f/�a&/*f �p�$�D�����	|�#2���r�>���`�W��0�g��,�����=�7ܖ\#���(��.6��T���BV�k?�_$�$�a��d���z�Y�У�H�ni�W�.���OD�A@gΔ�305^��Q켐ݣ4�S�����ݏ���� ��	&LmLt�?+��W#�F�O���p('}}��M�S�uN2=����b2�*���[�7l�9��+�b����P$�������zլ���J��mP+����-]^�es���j�jI�}ř2A�ALź��i&C`��4�if0����5�>n���ɬ���'���l��I��/�Rd�U�i�v-�Fl�Vw�ZH�v��� v��V�ʹ�<��MS��x'��0B����>,]���o�Wr�}���U(�i�喇b��dSwb=���`���A��Izb*##�c�`(�xu6)k�����=`;8��9��������b��҆��3W�@��w��b�|����3c�A�˒�&�ɳmY����#�χ�U��/�n�p�R�@G�A�߇�u��T�TW�[Դu�B���� ����xL����9����I�atB h��D�1�z�=���cj{�����H�ĴCNb�����Z-�L��HH=�U_�\�F�-���ig����%�x�B����E��G��Okl伃B�b"����K�H��m}5�%X�H`6B$:��dJ���� �z`~�s����.�5%�Ӎ�x\`Wf�c@ C�O.�m��c"�nV���^�=����Ew�؉�G]��c`�(�E'/��!���DQ���B>2�#w諱A�}*�R�D@M��<�59��	R�H%��x�"$U�M�#��U�2�<m��ϖ�,���UF�Fsh�5��_��J�C�PfxD3g��(�u5�������t��]�-?:i�'��u�,i՗]t]�L���!�3���C�-D���/�GLK76�G�A�i//wH��Ӈ-�4��U���bm	O�i	�U�H+�,=�YM�y����e<�G���,��5��b@ܜ6��e{�����d1JhV����Ļgݝ�18���"�޷q�8A~"�Õqr��,V�ro�B$\�W�$h�#HyI���<�!�.�L(�J��π8�z����uy�d � � �2w3dO1%��K�:�Ɗk���D��*RM��E���<��?�_Lߖ,��h`c����m9"�t��f���ؑd|�Ի-:oBM�Ai|�ׯ]�pvj��X�W�&W0>�x�W�Ip�Q��>�1 K�h��&��+W� ��̥��[8�:��vm�R��aY��֟���j[ $���H���
��� ����;�.|��� �O�x�NT�@J�N���`	��g-�����2�O���	ݾW�|���H�c�f}!8�~Hԋ��{䂙'�*�(pK�`�����މ�t���-J���o��Xh��?"j���d��LVƏ#��CI#T&���}�YL�aM�\`�",�8=��@A8��S��y����45h������ш[�K�3��b�s
�jvlWs�ͬ�w�j�Ĕ 8n� ������)"��z���Z�fL��mK�9K_c�*�R7����p��88��� ��2��`z�(~&��+��;��%d��z�#��4�|��;Fr.�Q��;���n�}��x<6���S2�� �c���L�:-@-^��2_�)nJ[��DU/�,�?Ɠ������VB���0�К�b��a,����D��U�N|;��J's*����ڡC�֓��AIⷁz��G�?�}>;�U�Z��x�F��]���oYr���=ma���H�v?��<�q/~��������d夺�ݤ-`�Y�vgʷ
�[�B:����g�/n���GA�?ێN�b2��&S���y_1�;9��J��X��?� ��5?u�m����e���jr�q=l�xbO_ 8���N�G�]Yt�0�P��U(AoQ�sn�/�Ӣ�P�>f��ٟj����ae�lQ<�S���Ic�xqe�L���|�6x�8�ց�ϛ;!@X�Huԗ��N�'l2�|��Hz: ��yR�B�н��+�i쓯 	H��H*z��8N�6ELn��d�Č7�U�"9_��>q�o��`���B� Q;� ��� �+0��U�n6�MQ�N��c9�����Gʲ�c-�!�n�Χ��*Z{"Y�H[^+�\ꏵ g8us�ӏw <��>[b�py��dP�yrw���{3*��G�C�{�OD/	of�V�c��K�f��⟊�ř��b)�u�j7���� �˒�S��-Mt�H(G���=L��!9�ȹ�<z��?�w���sP�M�t�j}����)K�É�>�H�c�v"=Y�a�KX�R'6������rV\'��N��qw>}	cjP�#�IxL:����k�>�CHņÁ�k�~�ˈd���V��C����yB�Z�֦�;ri}{�.�38���f�=TB�A6��Vj �E$���
��$�:�y'&�W��R�
U��l���>��p��S�zV�P�:ӜЦ�e_L+"Z�˨5���uy�2�Ex�xG��P5���HM�l<�u�C2�o���ңb�w0�/4a
HC�q�0��r�!f��^JV]m�l�1J���m�D���gB:N�j��%�J6(=w���&���],ǎ�
��X��I'�ߑ&�P ���a0��^��ܯ���p#���Z��s�{?������sc���i7˜|�ৗ!�L��BSb,��s?��±[���e�8CA=���"fVY��}t̒�������⷗bq����Y��n�35�(����g�(e4�v��%��.e3;������s
��'�B�S�I�@�eV�e����d�����T�]��ά���O[e0n�v�籼܊9�S����
�? e�����<�|��Jts��`�J�2�u~U�\Z_�o�x��?y+���
���C;-�J�����$P����sI�W�-:NǼ��ݡ�s`I�L�����$���A�Y ���Cͅ��w�=��60�ٟ̿&���?��2��>jd)�LW!PKA��J���@
~��i���B�G&+�r(��t�ڢ���W�?��cY"��~U�Q>X�c��V[ �� ���8�$k|`P�6}li�#��\��\?C!�m��y��b{QY�du�#v����
s�����o��aF.� oj{8d���'ol���Pf]=p�^���v����ݝ=Bx��_|}w�x�~
ށĥ�4�69$*�|�x8��$raօ�w�� �TZ����:"�˜`JLy?yJfM��W:���[�̓�n�^�gt�%��
��͖�.)	��5ֻ'#�.Q����Aryviޔ~ZU�����E�=���gcvl�c�k�0o~ʋ9��4��)��$銆�vm�\�R�B��BW��u��[�X�:��1F�����xd��$
Ed�s|,9w|@�9l����Ŷ��Q�61���P� y��m8{��/a�v_%��d�� $Q���R���d�RP�=17�Nە�Q/�����/6�~��v�v��G�m�_*�'v��d�l��O[�VS>���o�z��zJ�w���^PQ-�rII���� h��I���E�k�A�4<Q�2��~'�|�H�+�P%�4�����&��4�;�Z����l���\����;Jތ����)�n�BM�����<p�R{\�����%F���Pf��������W	z���D�H(���-vRϐ$�F��|8���:�ooHm��b�	��Q.C�B�R�gL�N5�ED$��������f`���?���Y��g��^@��Ո^ɣ&����U7�:T�}t./P�|�� ~�F�|�$𞳺�ٖߠ��F�$\�WQHg�G��R��?Z�\��!ݗ������hY` xDQ���%k<���ur�8�"^�R��p�*,nj
���=d�L����"<�6�ݓt/�:�v�jx�?�}V�y`(��!��AKY9�a%���ur�/-��$�X����^���EoVx�y�5?�d�8X��=�"|�r��\©��w-�����ā��sh$��(5S#��O��F��g�5F�'kj��*����:��g�u���!\e��x�'l����
��c�8�_$�C[��"��B�J�+xƵc�}�7��؇�� Z1p$��d;䒋:=\�4Q��m�R|���a��R�o����ج�7mh**�e���tF%X$��°X�3��P1��x������I�B��̨���͂6��jV�M��Y�̟m��/�D��	Z1]]�Qe��A�(,��S��"ҋ�����y�h�P����-[�P}�s�i�\�����3�M����|��$�o.�y",�L�L]���z�.�_ak�|�� �w5�լ��Az�?�L��l�&m���6��;������#�Yd��lb����|���<�o��=#܀6=={b��]a���B���p�����hz[;�����Y�C	��/��s� j ���β��w�M+îHivi=��ut��Dq,!r��dɥ^V���Z2<�S��=�]�Op�0�/q���C��D�2Ϝ�J����:$$'0G�q����NU��E���ٛ!�x�p�_g�,O�X�g�t��D�5�'��8J�U9J ��ܶ������~�9�JL7O�,P���sYf�h����.q%?g�s�t��Z�|9g��u��N�G�්�����J*��B��%�+!�K��݂#5A����A�m��8c�|�j{��u�h3	Z�i�W����ɲ���m�b�p�X�o/���{�X��j�d�wg�KOW<T��h���ȫ&x�c���)�}�S�D2�k%nYY�:��5��	������)�.8�d�h���<��o�/{`}�"�0��oR{��<��k{E�FCX���`8^��� �Ib/7�hH�8ھ��A��}��A����������p�A�]ڏ��[���[kȊ��MR���@�E
{=X�b��:��ҿðqV��阊Ԑ�8N��
(�RA��nh��pvi�=��y�������`eס���P�Q����!ӂnT�l�{a'��{��k����R���x����$�"s�ѭ:N��UٸDh*�`��@ʞ)�k�)%�@O҇D0���Ao*��eE�`��L�Ԣ����KV.�{���h��r�ǣ/�K�o$i��"������l׬K��AP�poG�Q@�a�w�=<���c���ߔuxq�U���Fn��̕�i����ħ�Q�8F��	�B����AdƵ����AL�q��@\�G@[f�°�K��l��mzQ=��{�gh�5��"1��@{��/��yC���Hq%6�x����~�I��!ԑSţ)�m;�i��FSJ��$p��2
6�x���k2��|�i�'?������/>��� �7<����0� ����E��O"ƹ��U���t���9>0�|����\�Q4��#΄�����yz�΁[��{ R��II�c�=�P�*h����
)�tđ��4	|�=��� ��j)�+v?`��<e �5Jܷg��d;�Ĉ9�G)�W�����H$,�%�*F�,�V���X���
�c�n[	�bI��{��#����x�%����;U�y�N�>�#�\B�x�V��7��9������������ݨ�v3m��������p��֛ׯ�����ڌ`ESM�w�� �Mr+���k�3�ׂ��J\���ֺ󿔋�jDPf��m��Y�����7T�Y�H#e*Q�}��Q��?�~M������"zCt����הf��?�vA��y7� "��������69�#2�.��PzH$I�ց= ��/Es��g��'��5�����?i��r��Y�-8�z+^�3�zl�!���1�+<0O���� ��*�*Se�3�hĕ��R�f\�)��#����mˠBPQ����PE1�� JhxI�k�Dk{1�W��]ݔ�~�U�y�p�I�%��M܋�����d^ɡῡ��f��f/'�7�mmRQ����^����]��Q����ˆ2.���qcnq��H�8����ڪ����Λ>���֊vM7Z;��aG��2�_�hV��d����:�T��/aA�v�[��@���c�G_'����#��S�@خr��ot]����I�XlxVHYEB    fa00     cf0^m?�IT�#��1#`�2�:x��,Nf���"1�}�>?-�>�=Q>�u�E,���/��蒖���L8�r� M��fϏ�X?��H��r�p�5�~CMV�"�J�'��� � ͱ�K�s��*�[��L�P�������c����X��i��Z�#��\�*�~Lc<nq��C,0��)���T�G�w�̶�1�y6Gh0b2.�>��3�$��1!��#��|mm-��k���T�`�
Xz�y�`N��N:��%��CL �������	Bw����I��'���/V[b�JWns������`�D�ƫ��^��Q}��b4�6��HL�0#ms!Z7B��#c@��[N;$�Zn}g���aM:�&��[� ʾ����Hj�=Y���cQD�� $s �zi�d|tV0��^�����w7en&�<�uZ�FA��9�����O0;	�\|0ݺ�n��=xV��S��(/�rqV�.�H�iyFo���dM�[!(jnf�����1��.6s��ȑ	Wf���a�՚�|5Uz����_*�a�'�����O����Sϲ���*^8��?R�UTB\�Immq^����),��<<[��f�s��tȼ/`�	���YY����t�'�C�:7!|�򍛞LAk��1EKZ�P����# �q�MՔ�Ɨ�<�6����yk�`3��-���|�jw�g�`�|�u�keİ�����8�e2�d�'A��j�3��h��� �4p�&�<5�Gt_���'��Y�
��U�$Rr��A;8 ���6��6��I^���	��0�rdQ%45�z�J�Z;jT ,������uX-��Q�Ohl�M-��Q���kg]���G��%�Y;mW�l���0��;���1j3��������7�$���%X��|c�d��:W�"��R�B�BP��q��|�إ)�%���>�F�xy�=;G�+�?�&tAf�(P,'�u�
}B����Đ�r�x�xF�x��+\3H�b�����C!��hE�T�-h���@*�`\�,.��V���b�\9��P��r�(Ou3�l���=���019~c��QI�8��]�V��l��*G�����sd ��X/�!��e���?��|n���B�ؤ����#l�O�Ș��LY����@G؁~�M)}80���u��}���یi�y�@�ߒ>�`�	~�^I�aU��Ze�\���ݼ+3��Kh�6Rl�Ե��okF���ۃHs=�Nz�(�;_�穖Ʈ3��
F����Ix]��"�+Z����J�mO�2�^�``��n�\tW��q��4m��Y,)��IWt)�P����I��im��l`����=y*b��q��n��2Z�Chn�r��G���.�w�@ڎ�$�Wt�T��"���5{+�E�>�^rOl��Z�«�w5�L\:L3�5�$_%�-�5 ��4�H_��4����zL9�M�Bw�ķ�_R=R�2���3���O���F8�LBs­�Wᒿu�����F�)�I�����V�C�U�q4�Q݁Y#�<�� �v�� �~%�ZJ�ߋ��~�L|�^�_n��K+��3�IJb�\������5���������h*U���B�.;���,�g�n��TX�*�S	.�fa ����2�k�hP��I������C+���Ju�
�w�^-�ׯ[1�j�60ÿ��g�
/�@��؁�i�1�)8��Ҥ�����P_�i�rʨ		1��@iP�y�Uc�����V������$���B��LT�HC�[�C	3�ml�kf
�6�o�Q�P�-E�*���3��9ȩn�~6Ʋ����i'L���P�o#B�>���9F_�("GbZ�A&l�W�S)l������"�	�Pc���Ό��@qj����,��&�\�+��n|�֗d�i�M�z�3�V�ܴ�#z��g���M	~Y2�l�%<�0��å^�`���q���^,f�����5�Q֕bj�Zj�_��*����p��|��VP��K�ޚ�����W����g�z 6YY�΋�1OA�m�ʅ��i���~w�ً/[�D�ʳc+�X/�]�)�F���ˣ�Mwd��[m	=����b���7Z�Db���ҟ�\11���b��;E�� /�ד>��5�#xʴ�ݕ���ų.e���Q\�j�#�����~��Ͽ�+u0��ki�9kK��Qi s'<�)L��<��C�ٵ�͕h���P(06p$�Z��O���_�8ʩ��)N�k7j�$j27�Zw4B�V#c~#N��/�w^�7�+ϟ��v���đ����	��Ў*��:!�KQxh�-k���/�h��@���h�n
�% ��琺ҥB֛�R�-�B!�/��bCv�^��[��~�������1"C�up��/�WÏ= .L��b0�YW�H�,,��?�B�[�~lr�&�"Gu�U+���,�rp�y��9\!������Fa/ס⟄v	 �&=�I���yY����f�$?�ź:��� �ۡ�J���ҍ��R&+��xr�wi\pQ-3![�%H�Ľ�r��g�~Zٻ���D�a����`2�}*���+�`�B�`K���Я���A)��cRm��,�@a5��A��Z7q�+<s[y��,y�)���p�b���iu��j`���Hҳ޳x���)��(J�guʰ� �(�#�Wb(�#�����[q�G��]�]_�SsZл����Ά`�s4��2P��Eq��o����4���9r�������v��qKB
���c�x������
��(/ހ�y'6��t��mК.��od�S������b�t��f�ɸ�ըi�1�$q`��R/�5��$�Y�Cv��-f������*���s�Nz��8	'��E[*Ѳ��O���PX��6�'�+z�f��͙��nu��K���{��>�(x�i��N"3�E�?X��7�5�xp������,P�=P��Gu���5 :��� �f*l��j�p0��	T��fY��y���r�V�m0�2A
*]��ã��
��WY7p&}�,}����gW�	s`u:�y�_3W�����?�j���z��	iFٿ����2�ƽI�_f[����x!�ȶ2y�'2z�dE�k���p03�,R�.�Fώ`�q��9���V&��=��0Ǐ'&�T��$���u*wjM��A�A�tkw6k��u ì"{�%1Y�>��h�\Vѽ�cF��F��D�
��6H4����F�l��p%����h��O���7O�8XlxVHYEB    3996     4e0p%zX>��99N�"��s=�d�f��	��������\��9��c�w��	��}*����ۄ/PK��𩜩|>���6p���;�\����=��BoQ�;��p�	�8�g+���3��S��}({�w=̼�HA��W����K�KH?)���@J�N�I��n<_2�IU�J�5|2��NB]k�ڀ�
Z�F(� Y��;�q�ܿ�8����Z��K�z���lq���RD4���BD+��ct��S�v�)�d�w�u�.64�GaK�yb�����L7� �F�-"���O�>q�I����`~L�h9���:�$�bVMB/��ؕ:Ž@�fB�Cu�,Sf2>e♊��/愋���fI�;.FF��������+�u��3�F:�:ŭ��{뛿gN�[� dQ�ׇc[?�b����g��#b�M��ʟ^<�	P����XtYa�hR\�1���Z��:�s>���nxsO��@gN¹�<S>S��&]g�v<Q��h]�g�5����Q�*���4�"�|��t`�����h�t'7Y�����msMJ3Z}� ��1ʋ|�ML�	z��{�!��3�!	��D��X���~�F4��~-���G��wг���d`T��� �[�(��"��D��4-�R#�
�ڟӮ���Zg�M���,���6�Ey�Eu�4:3�#�h���.�<x�:�ulP�%5O�`	�=u-i7���%V�
�k�e�1�^��E���6@r�@��,���tV}��(Qp=i���pj�|�V��]�����1R��=���H�Q��g�"�)���r浾������F�$���3XB���F�%�}�����X�<��������l~�HΤ��z��Kqh� h�V4�P�����ͬ�F�}�zf}�&������98,fs�xݖ�pDj���x5��Tʇ�^m�&7�]�ȱD�yZ�$ʞ̾:Bɰ1�AvP�t?g
�uę���N1y�fƀ��b��N �J�ڂ� ݞ�t�Gǁc��G?@av�����Ң���r��7=1�S=R�K�&ֵ�g�]�{��={��Z�������)cz4�w�Ȩߛ�*�I+]�Gf�zQ1~Ր��۬�S�N��w�g>��n9���\�;�nμJ+H;�f�����"������i8���o7%`����D]�E��u>Z[@ ��`���*��q��`f�vh�����I^���]�:�V