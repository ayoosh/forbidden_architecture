XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e7�d��P��O���7:qА8H�TA�������</�=W!V2�����Z
5����!����i鞣�n�M��l*�"%%�I��ADggp���]4���7�Թ�����k�}Q�͜�j�%d�Z׀����1�N�]�Eټ
�(���av��M��MT��t�~P2L#���;��T���.q��m���tXE��1RD�ɭ��I���s�юf�S��*�wH9��S9�BiA��$�bMk�����/�x|�"�/������H���e5]A�c��ڒ�@��㲴<��bQ$yD�>��1ģ�uO�Y��a�FU,)"a/UO� m�j�Z0�fÆ������z�?��P���[��,؟~�A��Vm���)����1�}��	���y���g��[HQ�QWv�����a� ���;�����bz�x��O�N��沣Hj����]~�9I�7�	!1/��4N�A�����Ψ�K>�� �ߕ��ڒUM�-9��g��L�T�`��PeHS�mcN��rn)�H��� �	A4�H�D��pQ-�N:r_��w���
����/:U݄���D�`F
J/b�N�!PfL�({Z��-N�k�{�i૥��5!�Y;�3��a���䪁�����L2�Uy'vs�N�|�`g��ׅ�w��7��'�yp��f�b �Ȝ�J���
�:�@'���I�l_���h�6�7E�y�k��b-�Z��<��t.j�3�N��NW�5����OXlxVHYEB    fa00    28c0e�o!�p=�x�J�B�A�咵�:�P�.�k�DL�Wp9��N�4"��y�`���?��u�����an�|�9��NYe�. �6��o�����|�"��l@.q�c�'�jJ�[�pE5��9�O�a���%R��ڞ=h�F���>�wb[�1�����̻���͛��wI�I�h�72oh@Q�&T�Z�?*��0�7%��E����U	�m�Mt��i��قs�^�*TYmu�)�Ɏ
��KQ`�$C8j$\~��4Z�(&S������-��f��}D1\:�)Z,�����x\\�ru;[I�*	2�!��ׁ��<�yg_,�/�2��*61�<�^+U�]�;��W� 5��]�_�8E�p.�#�1�k�lOaļ{%��a����]/��6�>_�*�φH�>�&�&ނ�V9�� �|-�7=���8p����^�ͼ~6gJ(:�%��n� �sb [d�X&�0�ޏ�o�?���(�q��,��(���K�&�2{��[��MWA�ޑ�F��Aq�e��d]�eᲟ�R�I���p�w!�l4e���3s��ȿ�SA*�7����:Ŭ��ˉBT�<��w�g�H�݋计Jy	N^`�XwB�����*�4��t��ʷ`�Kk���0�!�X�5�+�z��0�;�{�ǟ��\=��u�<h�c��
��c+r�<&������j�M����%��	�G&�5mA7�����j��J]< �/��\n����W�/R%Xw�X�I��?1@@��*M��_e�e$+��y�.�29/��A1��.��F��� <׆�$���R��o�Z�:��&�$�:�*�9/�G}��9O�dz�_�C�-Y��AUn1
��ד�D��Y�c5̟�m�m]���I8Է,Rx�ݳ�5�X/}���p��:z�~LXp��r�`4�Eg]+��}:Z�������g�s�Off;��M�7��ډ�@w���e��o�t `A	��1����!�nM/m�B��,T�\��R�ڗ���&�9�^ﻓ����+���x�C#5jx}���V��E�t�j�����i�̈1�-֒����N��U��{:�Z4�)w�~�����GY5���n.��i1W�`yKYI���y��fEN�� �KPvz�0C?��B-�����]G S�Y�C05�]_�}ǥ��i;�E<6��}�6�SR��<0��<���Έ���H�C�0�r�;�M�n���X�wB�����4݊8Kݦfzҵ��Ȫ+�y'�:�a�=�JB�P ���JB'g����t�5���B¯ߡ�X��ޱ�Û��L+��W��97U-�+�A�T�����0��2��é���uІ���1��	&w_^�$E�[��$P&��k�X�~��MZ*�3K>�����k�������rQ�Z������r1y�N���>��R�j���ݣ�r�A&qj?{v�IQ���ڇ~�1��.�|�D0ĻS��gbD��G������2��2��aFab+r���ܴy�X0�`�m@%��1FT� ��î^d��:c��I1�
r'�b"���-$!Qk� ��K���5�j4����"Ycf����C�P匸��wN�CӼ��z%/Q(�f�c��q_|���E�W�)��Em3UJ�_K��Y�����ޑR@�	d��2YE; �8�'eg�/X����)�]��1)&R()�#�7%��D�u9����/R~� �H�"K��Y���j�w�8nIj�{9s%�����)"(W(���꬇^4��md�5	�ӥ����Z�PN!�aN�NA�Z2=�o��dǎ��5�Qn�eC�x=�5+
��s�f��9�n���E��[��C�y��~�67	ܯf�gӏ[	3 �v"�L��\���Ǚ��/Y�ʣR���O3�<H��YK�g��~� ���ib4�x�5lt�
M��O�`b�m ���GZ�}U�oǂ!fgr'r�q{	�9�<�NI\�k�F����g��NA��w����gT��fyS~gGw���7B
Hb��7����½�S؇[1K�
� 
�=���y���{���L���N��5��UR����>�/��}�d�۽9���}��M��p���vn	D��r"�҈�Nl�����C\��<m�b[#fF�^��2g?|�l8I%(�u��B�Н��ܜl��*V�TR I����7s���6~� 4ӕP�ɶ����E�rX$�>4yV�_�e�B-8�mA�J�S��2,Ng�QՉ�����2��#VM�5v/��BC�W��=Jds[��ڗ��;��"�xjv��%�vIK����x���@��yy���P���~� 1��G�=E�'d2�(x�(z.�j�)�N��V�;"]�i���:�����4�xv�O�*%G�9��)�����qro�t$�IܸRq��;v\���:���ۇK�I"�x������L���H�HC�\��Zja\� 1O�5����>X`���!��|v㨨�vV�=R���������b$@S���;O���ԝ�i��2���w�&|G}7����G�2��C��xU~�9�[4;(%��g��l֩�!=�d]��|Bx�2ZAC����ꩡ�G��P�rDK��M^��	l�h;���sґm��������Ԙ����8w�����(ys����^Q�;�d���C�]A�R��x^��
_�ZBtƝ��7����W�aeg,o���*��c0���!���{��ʇ>�+ �s��f.`�- qXDG�+�m��6�'%�\�������}2ʡQe�o U���
T�:�#�ѡӋ&��:�ϼ�@tH���L�A*�{L3�֙��-������� !RqL1.ߏ��F���sF�%�/_�jۛU#Q;`C����V�:�f�j-w�N~�� Z�yL��u�Ch�Ҽ�*�/��Nⴟc/E�!!��}�^ �\;L��GvSJX* ��J���_P<O�O�U,��uZj� $�/"�\G5�tN�8�_�d�\t�Hw�\�AC����Z�M�Z�0u5/�T@��������@q%�{���[�F ��?}��4����Ƥ�ۊ����R�|9��k�r�b$�U�����.�ܤ_�6f\��E�� �4�K^[i4x�9X�Q5�Mk��%H$̹�6	]]WD���Y�q
�ؽ�����W�N�V{n+^E |ז��#]J�K�qxV��<9$��d	�:D5��,��QL�����Yq�ǘ�]�x炱Yn�CD��!
��!��;�j�q��1�I%x5�E4����Nt>���<Q�,[e"J�� }w�J���*���Z)ۭ�i�n����{8�;��������D����+Jበ=q�j�N$�qT���
Xg�E�G���b3	�Bx��K3�E{rN�.L%r��P�D]����5��7F�ǣ	�Ꞣ���� Mt>�L�("#Y�*`�0�eYy���%v�g�J({�Y���ɴ��VoΞ3�Y{��3�
�_�7Ἡ��W��^iF��,���w��c��%��[�*�Z�㔀+*���%�2F"�s�p �W�����c�h1��P��A���\(N��H�A/)��0#��b���e�a�3�$V���r.+{v�X��ѷ�s�2#�C^�0z�2 ���������L��aO^ҕ.��R�;�i�����Aku��[�e}�rƄ�H��㳴M(����UA�dC1]�2�I �WOs�5n��6V����m�cW���ͦ��o��:��|�	z"�lשV�2��z���z��� U���2q�� Z ��	$�����7����o��T�%!����ҽ��0�&���Xn& O�ʵ�ք�D��#��	O���j�3Jm-s�]���P��*�!a^ec��������U(=~ū#��nƳI�����[/��M�Y��b�<������#|*��s�`c���r�S@�J���W}jf�4Ӑ�C*eO�x�"S�;r�N��;U�{�H�K�>?���wިBdo����J Fz�j�dF��/v�Y��R�7YV)���5�fW�!�?���H3��]��(�r��kp��"!��s�-�b�h/��f�J,Я�o6�ϐK���p�^i��0X��1!4j2r鵆�����:/EI����SS�]��Z`Ė��m���#7\<!LHj�ǵ؅�j�ԫ���ˑ�E��*z��[�}���r��p4�O��6��i!�F�\�{]k_���4�����0��'h��͸������Y��P�~����AM�e@�L�v`J����=��o��}?!~�g�Q�c<}|g�O߆^���@C����w� Z~�]�<�[F��\��;���?F��	u�wm���K急���AK2U�y���$�����)�!\|[͊�k4rq����T��� �?N�؉׈4<]������m����}�d�B�U�	��������U�f;�x��C�Цڴ���~�WH-P�oܤ�T)�����gՌf����W�$�_�^�eǙ+Ԟ����Ty����[�����ڥF	#�>�j�C;q��/c6��+"�d]��Cn���W��42�r)]�9��J�R����G���"ыȪ�A�s�zw�k|7Y����Ȍ{�C�N �>���TX�o��3�61I���Fcy�7��z~�������Eξ����ϝ_�->����R�.�xJϵYW!��Y`C*S�����;um�JH��."�04;�j����dH��{�ZP�2����)��c���f��U(�7aW!��,��-���}�"ñ��M�<K�@��[�5*s����X3��!O�L�5���qU�QViQȣe���]������
��|n��c0�r�l.�Z�O|rb[5�F�*턂a��<^�Xf7F�C�T3��cd��W�yV��[����<j,�3����Ó][�/Ru�5�B�n�U-Z�٢�£�t��#-�&�n-�d��'���qb�崷����YN%�,"�3y=b�8 �l6s����Lk��ik�u��'�2j�GFŽ��zޛU��[�ss�e㥭��Y�J���}i�2L88fUN��΀�G�U'����㑣_D��5��4b6�KL�ͬ����	L��D���.q�o�gXvA�Pn&O �_�TZ6Pm˒&Y#*�5�w��:e��&P�"a�"� �'�NO�b���f@]x;3��Cȑ�
���p���B��<x6��
�Ts�x%���£d�p��U|.��F=�ؒ���?�|��ae�=���\������I����V���q<&C�j�_�?J,�o;3+N���[����%ʥmS��� ����㶋������~cx��ytL�4�F$�*��K%�'����P�͔�����j�����gWe�;�g��:�Y�s� K̢u4: {a�����W�Рa:��^��4T3�i8�6�ʌv�#��m{o��11�Z�����s��-��ӏ��#Ȼ2�Tr�z.����@Vwbo�セ���Xš{���m*zU�K��fZ�Ց"��rh��we�`�3�	+=�zA��w�T#؝�Rr�iJf��[�͗�Ic/�����W����SDKI����κ+j�UP�d�Sn�l_�34����N��<O���}E�Z{�nV���;u�~�⨘Z�����垆���~I��w������*�N?��/3X�P�+;�gV�]���g3�D�-)�t���b���v,]CX2w�>��_��:{��&��[�=M�ͶM��Hb�� �D�k*v_����M��"��Z�U�g<��Mr!qBz�p�WR�G���4V��59�(�'^$:��� �yS̒Z3��pwلu�nRV�k��kH+EPmnz1����fک��0Ƹ�b�k�e��In�t\�V�e~-��!��N�K�8�eJ� �RE�X�}l�=���}�!�dSp�!����+z�}W.�ԸĦ������ѫ��8�Z�S���%��a9�Ea{�ו$�ZJu�V�`�(��₊q�75 �6����-���{��rn�5����@S���e�����M�#�s���3�s�RCS��x���p�s�.jho�3�`���ޓiK���ef�q�!Q�;	�U*2E9�ؽ����~Cd��e�y$�Q ����xH�dp������睤)�(����,�D����n\L9�1��J|V����h�4�Tm6�~d�쵱�{7"�G��EoS��%�"�VU�c!��ܦ��>���Or�!+�l����m�v�y&6P^��[���y�*�}Wuo�W)�����Y�,��,^H�:��2T���M�a�z/q� ��>��jK�eF2abW4�$�ϐ3���I��ΦRxX���l)���:�L:���V���A��]]�	�J�3�W<y�+�U���C\čA��8�}?m�= �W2��vb��_1?͡�G�i�+ե�!��[�.��Χ�̈́ҊS4t�52�!?i����+u)�lח�[�R�	�� ���N���D�ҙ��rb����L0��u,�Oլ�r-��爳h2H�b�yW��9= G'�jԓr/EF�g'u*�l\��PeZp3��d�YHP����V�Tq�`�Y�ڝ��
Nħ������`Α��+cŶC�N!��W+��L�1��Ip$��^E<l��"�4�~��
`R���U���9�|���w��3S��M�`��( �z�,U����v�'�HZ��2`Hݮ�+��x�R�N9�=H���CW��R�bP��'����� �1�&�W����(OTX�ƽG�v�b�U;�(k'�(�U�X���1kR��A�r~�(hc�a0\�mr�k�lU��rH�r?$����5��p�kv��T<��5J4K����q�P����L^=�,���7�mS�$��/u�I��4����()ڑco$-��z4��2N����D�P�{�#��g�����){��6���*�nx6�r4b��^s|lp����]��j��*�S�$�P;�y���o>3zZ��R���H-H�aU���ь��׊��}{���P� M��Æ)%vl�Wȥ���}���'#�{�{���4�F|�$F�H��NA�~�k�/�y^ɤ� 8�N��H�(FoAǥ�`~�ZЀ	���mV�%�9���/gz��j����{J�WxӲ�����ސ$�N�U�|`�����5��E���m�վJWK�ʽ��=0��K���P�b:�>��q�O��d!HKT���L��P�RQ���ٛ��1����6�\�cOH�2w.�����L���������݀Q�eF��/b�o��&�����2�u�_�F��"�܍(�������]��sm|SY���Ӣ+q	L*J�8���񶀚.�r&�ҁС���w h$���[c��-�#��w��n|ف��Xt?1t�0p�8��.��SG��(DU-���+}��X���}���;�B4�^n}���P/��I���p�Q��gt���8�Z�A����2�����v��=���JL{�lh$�¨~���O��_ ��ps70�6���~(h�WQ{��/�[
��-�>�մ��x�T8�'A��G�1$��D�.��fM�k�{T��*�wf�Y�N5��HqU���$HNUr\�"�-u%�����g�!VDb`�*ni�h�Z�W�1�(��*tj_ੰr|�;\FB����6GL��V�WcR��3i��9��ʱ�^
d��)
�����6�N�{����	7쇍$�.e�#�2/�Y\�4��D/�������W������+_vC��ζ{E����1�lYW������z�6N�[����_��	�����vCs�5����^��h����G>4�uI��z�j�B�?"H�Xζ���Z�aB~9��: /�^|x���vrKT�n��l��<9�nӺ
�=Ō*�X���7z͋��f��Ӷ}�l�P.�$#.�.�.ERj��ʺ���07RU��^u����ז�����<O1Eofq]1 '�z����E5���8Ƭ���6�ѝRW�/�8��	oBĂ����0�i���)�|!�_�ʡC��?��~!���@�A�$�Еd`�Q���m�o��%Z�d�}�������<������oS��0	���T�b�yu�{�;���Ϧ�o�����;د��A&�Nfcy�I��{>���>���}�;g���Л.W���S��S��#O���L�Mv�6Y�@��4������ ��A���ϩ��M_��X�]�i��w�[�k;�L�9���҇�?�~�O��J�VOT/s1��O���"
(���7�A�*<�n9��.6)@��j�D�kg�֠{�o�i�f�Q3׀O.��>S.Q�����o,V{���5�S��)V&<�WR2�i��Mm�w-��٦�<�>a}�F�Ĉ�'B�Pgl�J�9��x�?�LG�x�i�c ��Q��!�Z�~�r%D�vc�8	q��;80,���j0�(<�ȣA��29
(�y��L*g�3}�,IZ�s�$*Ns�������!)(>����i�ش�s���(\�(��I"u�KX��|�����ݼ21R�`�ʓ[�d^E��E4��Yq.N�h�A%�o�L�
��[�'��-��x�t��cw�)��%4W�セbIfט����O��ClB����)���px��+����{ռ�G�p�t���'}�ɖM6�ܐ���H/��'f�V��j{f�v�%Z�7Ѽ��ϕ������G!�[��ݾ�*��%�	�/��5�*�xN �������a��|�w�&³��o��N��u��{`�X�P��N��d��K�1�dJ��&�ϙW���7.Xd'�K�DsV�����Z���{=(����5#'�F>�0}�^�҄��Tt�J�}s�Ӊ�E��<�k�����W^��o(]�J|�i99�����SF�K��@E�J8#l�
d:~NQGk��6�u������	S|Ҫ���w}����B/�79�~Ddv��.W�و�ʅ����q�B<kðuz���b�U�Y�!n��}|X{%�-�.F���.#�L��s$�"#n�6D�ET�!˪ E?�������|��\?̅�/]AO���
o�)�m���}BV�H��?*t=�=�����[}���x1����Dgsa�s��Ό�� ����+!���������ˢ��U��K̳��
���g�[R!u@�1�Pb;H8F�P.j'I�ˑ���<�"�E��@�b��`rtR J���"� �u�����>�%��������9�D������
�W�I�0 O�	�#��ph�����	
*�B{�Y���Ov4������n(�!㴬�ݍ�o���H����G��{L�ޚ��C[?�3��P6���"���F`pU:��L��S1�-"�:��g�?߽)�%��+"�&����24�K� ��:8�ߚ{H�������,�0���ǧѢ�[}QP��ؕ\��oɵ���3��'�!qE'#�:��Y
�\h�T�%O�]h�|g<:_�Jp�o�f:U;|D�uU�+�
�C9�x�n����p�7�"�(4��IR�g���B�Bx�s�a��U��a!�4�q�l!�YLx���J��j	���r�Hj0(M�wF�ê�4�U�7!�<�:?��k@Ը�	�3�3��PZ�����m�޴oEA�	0
���bfv9���)��y�f��l4(�Yn4C��P��sԧǿQ"���r)�{ƽ��cؖU�5�ׇ�+4�z�tG�0תs؛�Z ���&�#�E����צK��t��?�
�$�\>	�������Z�|���3�9n]9�Yj��0E�;��t$��,-�@M���N�̒dG]I��|�����1C�tʙ���L�5���j�{����@�>h8�7��5��NO@�1s.��2k1�~���e­|�#r�=RJ�^690�����Ilӷ�'g�b_�"�g�Řz�>�ڟ�9�����@�(�|�u��{@
�
o^j������2j�f��.��O@
��]���U���keB���z�w{5�+C�s�����S���W3fg!��}V��)u��fW"�����,<��wŪ=}qoM !��_�u(۹E+n�d���Wp0�p��T�d�T<�`������_�.�-��I�%�����T��$��=���3x�Q|���2�y*X		G��@��	z^�%lXlxVHYEB     8ab     290&���.�Ii�:��ϱZL��ICǏν[8�����E���4�O��!d�|�������T��4=�#9b�[�}�HZ����ΥF���9rmj컗��ڞg��XSl��RxF�E�+F�w~{���/Q��S1
l�ZNن���1�y�_����~
Cb�l�!��?^��u���G4� ��MO�w�Lް�N�J�C^]�)��NM���n�����1�TKT�m`<yg^�~s���t�cyj0�fcz�`���%���a�A��=w�	*#O����i�>�Ӿs��~�L)�0w	���k#)���(ոR���Qggy%�痩�)r�R�[�E�%������k�ꗭ<&��˨�N��)��>���itE����?����s6��g4�D,e�Z��%��)����=an.m7"��
���L��bKY�)咃A�j�"���9��n:�-�\	���g���Y�q"(�V �̔b*�Pz�pJ;H�D��"���J����4�^ ,E�N�6�m�]���]����W��\���¸[D�c/�9>����"�a�^�Im����j:�W���Y���+����xʽ�Hl���Ǖ�Уx�
���´bw57�Luv9y���Z�ӕ