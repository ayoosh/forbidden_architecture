XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_�Y��+��}���b}�Uv��u�@io=o��PT�m��S�o%�*���=4��/2�x�QӐ!�9.��B��4M:��g1)�C��y���W]�tD��]�5���H���H12>�HB����d�.��_��a���z�q��y#�;vPb��!]�����"&��9޼� �8I���ڛZC�����,=JU��� ��+�@�H}g�D}p��T1;�;�D|$<d�y"������ʿeV;Y�f��:-�kgT�c�ٹظK�;U�ND4n)��H:�Q�0G�v��><�/�,��H��7�Z�1�K����-J"�2�kD����r����A�mʣ;{ؗ4�!�i/�ӥ��Lb�v��T����ۼ�`�ce�`�Zg�(n��B�6�K\=���1�|��ˇ����Xw�h��ׇ�rP޲���.|j�k$�g�nk��U�ۼ����)M�����"�0���a/b�S8�1�V�ܴ�`VD������0�(G�" ���<����5�< �����un������>�]��O�q�"�d���1v&%| ���
Bj��V��'��� О�<�'��O�C�I*��?0q��=o�_��x�;��:R����	I�cC��7@=|v	�-u_��:5��Ο�Ͳ2�aҒ5j3��^�*5�~|5��6
�g�]������W�ǜ�D��m~���(��'����Z[� F�����{���h+5�11v��I�)�Rì�Ƞo���XlxVHYEB    fa00    1950(n�V�NB}<�O�4söf�ڈ����`܉\���&c!���b�\Cևܰm�� �~�S��8�|�j�����1Z�������������b^%�O^g���ή7��a��5*Z^U?Ёr^1�/�ˀ��^��^Cb�����t� eH�^@A+�5i��H._n�"m/b�j��7�!�����b���?��{n��J�#Y?+;I���w�fU�Q�G�"���-|i��ņ#�c�}k����!̱�|�C�� �����C��V�ok�G��F�~F(,#iܝ�
�J���sD�V�	�r�x��	�� ��G
%I ��Z�ܚ�3�C�%��O��(�� T�ٞAp�Ѥ���ƨ7&��F1�Q�t����M
�4b�FD���+Y��rU�?J��J!���,v�\<I�T���~p�/O����Z�wQ%|$F>���L?U��34�y�v~���Q�B6vu��5Lq�0�n_K<wrI�t��X����&�}�L��Fg����D�b��?�[����h%'y|`^B�����Έ*��@)����ls�n	�Nl�K{k��r���%
X=k��[�탞�cO��d<�����T�� ��7�A�g^ %�عE�G!�^2����P���XW�6���ӥnH���M�5���j��K�|�=VG������43ff�Bj��hv
���dv��k���T�ej��6�u݋$n�
��Dъ���������)��;$DY�U������-2�\���A��B�ߡԤ�P���np�BI�b$�C2)� @����\|����$`�ǃP5��B�Ǎ\A;c��M6�2׊1B&D�Pn�����W��]hDH������wC�F��=1e4o�-[��!ڻa5��muqХ���6cw:�8C\��yZGRu���.k
��ˢ�(����Ov/�zR�;�Ѯ
ď�I�v2B�����^�HĜ4�O��Ah�����d���{0���k�r(�X��o�.㣷�`��d���ďi=o��Œ����f�����E�a�g�g1H��%�2<m#'����%��Rln�:�
�E��s�ʧ��}��/ðc��굶Ls�}���B\�>�
�R�F>��q�0��w�pl�3M�b
�
P!T��,���
���T�V�_���� �j���{Y �ӷA��D��Zu�:�w�V{.���G�9<����3�r���w&G�ca"6S搤P�*"o~���+���ף9L�8Lb�3�[L8���[��fܴ��*Kޙ�*jS�����,��>N;�^^U�M!���_$H{Pb��c"��ۘ��p�!,��H_��_f2sIV8�b~3�d�W����	��m����%��B�,�\��n���O��Z������ 2����%M;��A����J��u�;	X��As:���d1�M��U��䔖����[T��T�	
�dʮ��#/Ϸ�xٻ��븬�w7e��E#w�����Z�?�2��	�Y��?Կ� v��ǆ���3Яw@=R��_w�!�8���iz����'	���%u��?��9�*^N�V^k�@���1-���(�1�Ŀn̯-@재��JJ���(D��)t��@���Ӛ�g�JQ�0�u�8�^����*�*�1A�/�)���O7��E�����vYF��8�����o��d#��`ai �,]]��ӵ(:�޼)�)�{BnS�B�e��֎�ᖞ�0�^3��>���ܪ�@!��M����Qb�ZGǄ�4�A������I��T�w�䈺�U��!X�8���#6)���D�b�V�({��?H�ja](}�ZCH��k�9}����A�q��A9��6a�n^ժI=����ڽ��� �+v
=�l�*;� 1NK)$����zO�$4 �~�	ܨy0/KeN��)����[U�4 L��
C[C���Y:�ͮ�Ĺ�	rÔ�/Rʬ��<ϲ����1��'�F����ֺ�M.�(P�݌�3VO�� ��\x�i��,SFI���ژ���P���2�>E�mG����-c�v��D�J̌?���i�H+�."��t�txv�쀇:�0kdV~#�i�Y�������ԥ.er��eh wn����c���LEE�s�Tf;ӛ]�̠۬p����O�U�"K���@� %]�� �rw���L��<�Am	;�ۀ�n����Ǧ����N�D4i�Z�|Z
Abf�|:��R�"�	��P-4H�9����%�.�y�0��zS�z��6W~�z�&�R #�u�*���јH�������ZN�`�	GD{1�s�[46L���e�y��&{-�Ʋr��"�D{�)�J�DX�"Gf��A�ϖ��p<��������U��W��"[wT3�g�L��6�ɺ�}�m
m\]/�~�������B�3���H�<,��H�V�s6J;ts�g�+��h`�z2$B5��HԏR�(�#=���\��ָնT�'���Z��yإ]�k{�"����"`�b|iuOm����N"�����|.�N�W�Vyf�5�Ϯ?
�X�o7#ι�"ɯ�~y���R�w��%i���;s���~��R.���"�����`9C�/%�������-���W���ۗ4��('��u�$/�5n����E�q���"9��%��\r'���.MG�.
V�_{"?-����`�U�|��{
nJO�����=�&������RzTC/������$��$;�`��a��8�a=��|����'V�pv�/&Y�s	�P��fj(w~�@n��0CA���A^o4�
_B�G�UX����N���U�$����z]>�1��Q;D��
B�HQ��ZC�<1�e1L��RBo�o�9%���,)�L\���F5�����d/�Ώk�&�W��<�G��Me6��4�>���A�4ʨg}`���*-W�D�j(�ʽ�DFh(��!9WJ�-�qy��x�6��i�+q�H���ӵa�i�� �O̼q"%6�g�?5���f��������"W�ǩ��E����^|n�z�����vd����N��B�	�Zg�|��~���Aݻ#B	T\~����/�$}�qd�F����ci�����*���$��4�dr[��?�yMmz?0�U���7�����Y[1/��и���'_jgT�&���2�����N"��2��>���1&���c$�����bQy�B�Y��`��8�>Q�^Ipb�%[c9h�uø�$��,���޿x��������G��r�!w��$,I��;$$���j�Mb>W	\�/�֩����#v��4�\�����EԆ�9�^�����y���UZq5P��%�7ʌ�]�\ljd��>�N|E.�Ү�2�BM[�:{��1����I)m�S%{"�6w�Ѭ�g<?j���y0�
h\� ��W��M�?ô2�z;n�U��]A��ĳĵ#�R|�����I�`���%d,�FJm('L�3C3E��|�eõ��B6C��+�.����	������s��ue]>a�O����lCC l�-et6��X��0�H�jt�}�dp4c�{n��P*�	e�[S�!4�ϱ���)������4]�O�#RL�Y�:3Z�\��ᢧ	���
��hn5y��3d�1P-6YFT;�n�������4���I���]QK���3�Eݺo	�)yX]����	`"���&�Й�]|X��yxwu!K�c�d��� W׎��&��4��}�Y�vs�3����c{����3Ȟʊ��_����������u��ݱ,?#� J���(��6���D`-��zuۄ,�(8�U�E�懽���A����yG��x�&N�FH�~A���H}����M h:,W!R�mvPh3�\ȉ�6x��\�x�}*|cSe>>4��1b�s�L:���8oF�o���H<;j��¶%�,�J����eg$V����˾w_S��\�ܩ�Q�]x�\!�Կ���#�
�g6�$�}h���!�L��uu�^&�PPS���$ �����A�J�>�5� j���`9�h�|�m�e�ݔN�-4�e�Rbt�E��	�s��is&�R��HD��PV@�� OU���ZXBf+�m�F�e;�y�v4�{��p����-��@�vј&�z%��\ʈ�c����t�4c�U[j?�j���Wa����S{au
�Rs)zG-�?%9���r�ؙ'! ?B�y�i>�f��P����q���NW��UH������O ���K탃_ac���)�q��WK�DR!���y;S�1CRY@�9L�t�(��?t�JF;���N� e���K�g�u���,$��9m7�̏3�2�������%�-���E�;3�cƨ�J��T0��c�5D���7ǟ��7B,��o�4xȞ�]�ue'ִ;�{Ly�OQ�	��Q�������i�a.��Ր�����=i�FJ���h�;KE����ѳ<�;�I��昈6_##)�BMH��#NN�`�i��֣�Y|�֜zy�t��Q-�:}i���W5}Co[��|��8����)m�I5��=[��� �L��l90�)m����JoVTث��߸��B(�3;f�c� bY��(�.t
a��Tj��:�f�3�"q~����c2�0�z��cz	���X �����G�<��cm����fN/�[�Z�����V��F�.\V�܁��_U|�pc�,���]���c��s�Ő�� =�������r��A���a�C#.̳'T~Y/�{��u�+7У4�6;�k���A�QU��(�[�L3��E��Dy1B�@g�����G���5��x���M8[L_�\:��%)� A���)؛��Ş����t��0�po�(��G	�T��8QW��v��I�`�?C �
rQcCֻ7���l+G�5�hC�#;����]v3� D��z�0W_�+��
����e���.����_x��Qe'��'��NBW"!�y��b	F�}�[�~��2��e;(��Hb+�w��D\%D�[K���@K�bX��,��hg��fL/�+54$Ay+.v�0�r��4����Hԯ'Y,��
.;�֯HL�H��ΑD�'K-d�n�����.�%����p[����~�ڠ�e���Y,X+h&�%OJ'����ԭ~#����2=���V�W���Gϝ
���R�I[��#� j���;ٳ��[W�0���X,��VR����ug��K�r��MȘ �v��4�/�ߠ��U�a��6͞���b����I7Q���NQjn�8����⽑��x!r홳`�-�j�}f'��}�o��P1u�sy�s��s�D�0
�x��s�ݲ
b��㯔�%�O'��yT��y�oT��g�(-��(=�c`�83ۧ��Na+u����t�?��0�U�_SW��R��Z1اɬ�N����2a��tD6�����i�<J*�����P�]�X��,��j3����}��ް)�\H�$�Ks�.A	EP�p={�J|��4Q��4���"Vx�D�a␮s.��=qN���7N���	�p.�*��؀bc��@�*2��_��c���d��w��P7.c�#�n꫁>M�����~{�h�q�.��uw|����A^h3�,+�L��oظ=�[�-���d�7��>�=����(�B|��źzi���6��E�#�K���y�3��z��(��az�������Ҍ�[�gʬve�PiC�~�8<EاV0�x>��_�S���]�B�k��ͽ�be�yvXyhUl����/�N�e1Y��,�Ե���M@��P�B3�ҽc>,Ԟm��sP�MmbT*P�>N���*{t��j' ���?��	W$�R>���`AB�d�}�DS�QP$�7]�r��o<6��ڣxU��Qӿ���������a�x^ߑ�b����W����Z|ԡ��2�cWĊ_�W���D�F�1�Q�H7��"_>�Y�#rӢ��F���S�M?�����O��0�-����}$�a�X�[c!�nql�>䊶��6'p4�k4�X���(�ƒ��z&:V�S�R�ADBc5�:�0��qF���nVF�`	C`?��8�ޞϪf`Z�k�1&�=�F�w������F��j2�3˒�<���;�[7�G,^�EEz$�n8�DЖ���i�߶�38ޓ!���׫�C���Kz��=���)�w���:[Gjh�FzI�`a/��b%���#Xy�RX�昄]����/�C}cG���X7S�%D�>���C�҉���,��X�0ݨ�䙘��Seمi���:����X��$�fB2Wؘ���Ys2&��.
Ă]4�a�Ţ�C�hDآй��`B�x��q��T���PG� 4|W�;�]XlxVHYEB    fa00     700�s����i=`4�6��_��z{#�^�q[B�a1j�����7�߂ 975@Z@�9����/���J�9�G�@�޿�D�v���Mi�{��A+9ȸ��5%$&K�����L��Rs1X9x����M]�]��G��I��)'R���sB�K����}��&��dȜ��昻��> Nu�ئM��{��W����AUz��!	��N}vH�j3\b�T��Ǌ�Ā����~Р����#i����S#�t���&1���WF�ES��ÍU ��9�h�oB�����b��
���:%jG�2�j��6�rX���]��M��+u����Wb��Ц$�����'1и�J��H���d_��iE��A�7j`y�����JY6�ĵ($XQ�x���1_�㾱鋘k	�>P�1.��kxK)}��%�.�=���F<�L���Q����C�B�Ө2rK���}Ը�)�mV�]���&�a=���Ꚃ]A�DPy����D��V�ԭ
�,%�	�zu���v=�����ݏ���� �~
�U�X�
�$�Cdi�VO���rYZ���-Ύ����!�����#-���J�����ݻ�p����7���2
�V6�T$q�I�$�%��w������}��sa&�jqW٨S�}�I�Y-�����̢O_+7AF�����C�U^e&'[t�$d���Ő)�(!śOP[hf�n����Z���}��S�W��A�l۟|�������Ο�>�6O~��J�7��XK������Ң��ǫSkW��r���~�w���qB�P�mMs-G`h�Wl���3����a�\�a��b�h��ѕdu�1����U�Uň�'�%{��/s����L�|B}Qp6R���~���<Y+�lV6�[H��!1PR���h{��A�y�т���۲訁�f�B�a�����xh�ϏK�?�=r����YDROR���e����R-U���7�Z��/�h5 ����qQ���� ��� � ������<����u8ˢ=U(�G>_�結�-PI��NkE,��,����*١��-�YI�{��Y�S'1S^?>z0	��%*��H|B�ҥ�>��g��ٕذ��L��N�*���t��@i�����"���$�,@EKZ�7`]N��X�1U����͡~BQ�B�E�_|��U�>�#l�L6ӌ(V":��r`�A�o�p��XM��zx����M8���m��a��c�-z����.����!l!�4���C�@׀�;4�V;���W��|d��8��������c&��t��?x�����)^Pd"<�m5���(��j����=�
�1�8��@k+�����.X0|
���--�|�o���s�9m|Ҋ1{%�;״*@@)V�I�5�t�!J��c�*D��J�l%�ʲz�>;���������'��w�"KRc�ZI%��~�.v�B���?P�.�D]������K�^v
D�k2�}c��@�R�t�Ȑ�$
k1@Q�d���&J<�
}~t��b�u{�g `���m��Rj�WG�rIk��U.m̷�9��&�EZ�Z���A��&c�DbZ�{�ߒl6�7 ��VxJ( 醜�4~������	n۫!����z��,発YN������S� 2��D�?�T5���ς�T��|��t���Q��O���֜�6��7�I�=�"������[|�L��}�q��D�+-��nu�eh-:��n[�_�`��y���z.5�@߸�t�C�Lsyչ��0��%�XlxVHYEB    77ef     a70�U�/�߇5o���n˕��*�ێ������\��1�� ȴ.`i�p�	��a4YO����Zٕf,��������dp+w�r��@�H�����vq?�v8�E����D$�K����W�=`[51�P�ärf>�����bZ��#u�y6�π5/l��ú�k$��n&�'-�W�ȶt(S<7���%RԪ�K�1�\���oB#�	鶕>��(�̝E�@Qk� Fo�/ir�
w��P�E���đviN��D��l����<xm��3�k��8���%�c>�3�I�^X�B,�G&�T����&���ȸU�j�=t,b*�&D�A��U��h��v	
�����4r�?�<V�WJ� �0�'���6&(nş���{��2�1�CZE�y���5�-g��s�?b)�]H�'��n��X�ro����4�a�W�b� ~��S�*a;���`�k��e0G�]~D�l�P�[繐J�kj��c��m|�8�|�6yP8�0Tsat�9f��՞�R--ffyL�~��{'s^^�{{��BY�ys��i�������H`L�娉�|EkǀJ?�M��I�\�����'�n;f�C�׈�^S W�o��"`�Q��=>���x��x9��\l�(����e6��|:��g�K��)=Vpp3������?h#[^��0�7ͶŃ�8����E&�#�FLZk7
�B��U�n���X�QԺ��\\�	���Ө�il����)@�,����>����7�����	��UM�l��0qB�9��K�SI)�c�<	؅u<<+��a2T���ԩ���'���*�̴Jgr���nBe3�EZ��ɜZ�~���7"���g��<��H~.�)��ϳdH�gj<k�?�/�^�:��J�I�<1��
x�3��
n��{Y�(��)Us��Z�G�ѹ&F�M֝na�:��P�T��Osd�yڌ�Z�[�7��S���t��O�Y�b���f�c��dK�i����5�v�������;����}��c��vF��v|�@�2�����a&�ch?h1�BI����'�ښE#A%��s	#V�A��9�_a?�ɾ��k#��} �rщ�#=����*Q�����7m��VKCy�=cR"+��u���.i��%$�u���?���A~�Uwĸ	8��%�����"���V6�բ���sJ���+X��Ng�&��Y9�i��nQ�&�h���j��g/b�:�J�;��s7����=.{����S{���9[��92�s���H[��ۀ���P���|��m��F���K�3F�`4�T�
����M0^=��s*r����N����LCc�/�Tlƫ �w�C����$���Og�6�ɨ��\
z;��+��/�uI�����C�A-Z��r�v�{:<��X1�6�y�����G��?�^���lg,�:��U�Շi���$&#�;]х_�~�)S�Q��\��'h���g�l�z>Ʈ�W"M��-	�(<�%���`:��Ynt�|
��v�xRN�!�q`���3K8Lr������W���M.�&����s3�<����?�bTq�L���}��3��3��f�;h���s]3&P��s�Kk�A�d^��p�P�)MŮ;�j��z^2���W=�E0<��Q@I�o�ݗ=��/2t����9R�ol�r��=�b�G���X"=H9�PM �wQ�����q^߂e�����g�r9\,e]��r> {�c`��$mRX�u��T'.�i �rr(�~�מ̜�b�+;r��ҕ�[���M�\����!�/�5(�$'�&H	��ihqmx��*<7ۣ~�SV���@�উ�C� �G�p�w��-��O�Is�Ψ���D5+�;;�8�z�̯�J��;S�धI$m��)1���e`��%gb4��t�ג�[C�����{Tm�ؚ�)D�/����(L�[�s�-V#��
�2�zaa�\�,�B.��(�C�満�\ﮑ�d6�'�w2^�r2�*�W�L^\�FƉ��Tъ
jZurs$haU��2T��kӀg�����g��d�q�������*�yv��s�ۼ��MEAYՒk�3���#
���a�@3:Lj<�Z��;�~�S�vXjU	�d9E{���g9�Ĉ;�M��X���#��X��<���G[~ط�}1�[xn����������_��'�8D�s��uޥ��Έt���np
f\�r�Η%��LF7�:�1���l�B�}�IBEHl፫��F�ʷO�LL�<� e�����=���zD�E��Ҹ��߈m�C�P>$)�Us	��IL6��?�bV�8%�sc����(M�*%��^���i��G(�ys�m��NEa=)(P�
(kD@�mj��_K~=���N�|�w#�$h�^)§�����?X�)f��!3@qx�!7���ΰ�[nߝ'6�"�Rf@y�����cV�f���01�P���I�An�n"հJH +�6�L���j���q�r=w��S��~6�X�Yr�������a$�=7(��%|�9���O�l����\�qʽ�nSBT���^�_���k����W9���4���y�`��Y���"V����TH �b�t}p]��_�9�5/s�[