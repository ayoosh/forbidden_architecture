XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W�۝�Uڗ]E�>^ON�t��'���M���2���+_�B��}��\��g���j���BU�Ai�FWrC�_һE�]�8T���,⦮���W�N������,v46�>�� ��)Z�i�9���%����'k�:�����EE2wk����x�׷ߘ�d}�i��c���`�2�(��C~&�</�6� f���C���Ĩq�ʏj��i�vj�� ��:�i�������Z<�x�=�i�zm¦Qg0cvY�f\~-���J_3��y�N�S"�+���g_�:7���ǌ�W=꽞�s����ƶ���vf���F��'��:A%0F#wd��*8�ҡhk�߿dlG�{�+X��E�d!v�������$b��yIn�6��Т�^�o�2����L�Z� a��%�z���#��<���[.��cG"�}�3���)�*H�u#����4|Y;�(x�G#�r՚� �ѡ�B�Ch��Gx�M�Q9a#]Vۏ.$���)����CQ�1z�w/�N�>���R�� q5�|������R��*Oţ'�t��9�� ���[��ND�������y��OY�Ml���ˢ��|���:������YL�?S	�u�i��,�
u�J�-�{�g>ε(:�bޙ�G9�e�z�" O��cvO����ܮ1h���)�t�%��>��ҏ����9=U�R�^�k��
-���z@5#m~�	��dKz��9����|6��,�u  �fJ�~����q%���XlxVHYEB    fa00    1790b�wU�*PY�6�ǵ�X��~��_�/�S#T���kc������	���M����PC�Ue����#�=
��-�j���]��A������xF��5�Nꛏ���,	Yu(��P*Bѱ�l�)���J(b�X�/r:�Q"[�:'Yڣp��h�$ ����f�q�����4�*s���"�������W;�
^��~H�QH��'�MǾ��"eI�~�
9�-�d��X�	GsCrq�$��䃀g�͑�{jG��zR�!����7�a:����Z��WT�f����T�į���ۍp �ԎF���.���T/�\�!����kt#�kn�{Ԟ�+���		`��ϋ
�&p��(l��M�ö�8�T}��γ���IԤ��J�9�ӑ���]�My�%����T.��K:�6^�*���Z�$�GPR���gBז��,3�r��WIB���,F�_a��C��U��Ti*C�gZ��Ϗ�M�?"/��U��ŞP��A��i��3Rh\G�R1/��y����d�ݢ^V��
k�|���'�콸���3��zf���믺�ү/%0��\)�y��5��\��S���~��?��<u_Gg�^���W�Xoo��7� �p�k��pb��L��Wd.�D���I.������m��Ň�v�gd����!��|�aD-��*��7��������f��t+��׶"hN�!;0n�U� I�N���Z����e8���:�
��3� P�{C��Tn4�3Dd�?�����,Ef@r"��8}����MG}��m�8a�������O��K�5ߏ��j�;;%�s��.-ٻ���kl��pK��ӭA\Qf��xݷ�Rj����C�+9)�h��8T�v���V�lRk��!�a�=,�
ߞԫ�R5gjNvQ=
�<	Gl��۴�x�k�ESP��7*�j���&*p����ޟt��ܞ�K��D88֠��f�]�ȶ:�ٛ�ڣ:�A.�z[�Ӄlq�����J~�j�1�s����o�Q��DV��Y���T�@YX�H�&��n�ܡf5T��Cqpǧi��(Ն��r9mL}
��: �cU�X �x��!��$���]n�#��T�� {8"Ѧ���������>��~����i��p�u�7���/6�,%�i5��o�����O���H=���(2�r��3���]ӹ�WQ����#.ӻ�����s]/��:���t)���4
�g6��%���s�Ψ���%A=!!~HC��v�C��S_�,FEͣrCD�C�DI/-Joq#��G���h�n�}!e�	A	G��6)t�_���7�lq�,4 b���9����¥`U�^��Z
�=�S����zL'˃2�e�q��iU��d ��q�W1�J��Zi��������{i��5T�d�t�-V%���y�0�Q�V�a^�0ݼ�����]�7�y�"�/'^2Oϴ#����Ʃ��K�*�އm���	�6�N´�;��E��4/'J����J�䰱����G�dу�1pZ��@��J:/��Ģg\}%
g�������ߦ��L�ց��l�Wmy��A\���}NpXb�ڡ�8�mģ���g;���
om@~��R%ã�n.���������>(ϒ���AA7�*�ܑ��YQ�*d��l����X"J�&�L��\Ez% �e�m�L3'j~� ���s>z�ǆ�U�N��!.Ï��"V���"��9)�LtF� ���AH�B��5�[�˴�Ө��8��TVA���H�<�����|S�"��<[���F�1���D����F�罣qШN(wj4��O�Hk�e�;���I$<�쎝kp��Cѩ�吋�����ܾ��`����r��^���9E*��kY'�PJg�J�Z<T�SB�k'�{A�8��L��/��������[No5D�U�֨ֆ����oy�� �������^]+g'��"[���R'|\Z�KZP8��|N����2:����|��#_�Yº�ԯ�]�60`�V���W��蚯߂�נ�H�|�'�	ؐ�X� re��`�a1Ͷ>���f�n�qi�l�_�_\^��]w1�F"�cr%�>O������d���5��������09\���-�t�a��<��9��թC��fu���`�z'�:�-����Ϥ�p0�ʑl��fe�[O-� �R?w{�����F�z1�����<�a{dk��.�bB�	������5�	؛;(��O�+�*\�ui�z�4e����Gs�����	n7��C[�l�k*��LZdr���18"���W�L8�k���0Nb}�u���� :�R��6��%f���yv�����-P�|m���\��J$���x�� p+~�M`��Z48ܿ�F��~�[*4'9,ʢ;9��>��'�N'��Jd%���j���{\��\"-�aJ3@oڹ�����3�{�wݩM�7&3L�z�SY�<U���j=���GOU	���s���,��z�����\�_�m}��I����ռ�:���<J"�U�\q�Egխ�+A'�}Ì��lq��Aۇ����~�9��!N7{;'��?�_�dD�v�҃[6�ߏ�n2�2��ɲ���1 �C��h� �*�pe��OW.8��q0���||�_���v<f[��*xyig�Mʂ�� ���d� �|��l�r$+�E��HwY�.���e�"�Z� ӻC;��'֠Xت,�1����/'�r�SZ��rD^�� �l*�)
Ge�BL�׉dnܑJ�uC�FH���Y�ޮ�����\z}��w�����K�>E���G�գ�4�����C�;�i�h�4��l+>z�5�9l�iH]��U���1�O�� �܋i1X�������qf�|��܂�?Q\���(aI�TͻY���7=���8K7{�:ܾ6sgb��Z
�`]�T$ە?�Z���>��/q����-���~}A#�ڷ9��XS�r��<���D���t��J�{O^:�zZ�u��6��{���DBYFK�P$̾�y���>]+�ܞ�b��~	�Y�Y;��$��B�H�e���,׆��3�����l"˛h�5�XI�zE�LC�m�D�O�y2Y�+�n���ӗ�W/���I(a�/�xn�k(h�T�p�>�i��e0EDK��Jd�y|j�Z�|ŭ�d3���j0�U����C����C�}׊��I� �҃��Z?�nhV��Y��7�&֥zY���>��)Qh��Z�L!,U���^��z����4��KX��z��Zjߡ���ԡ�7k:A�k9�:���į���\�0�5�'���X�.5�ՉJ^hWG��w}87&r�����cNYbi�~U�/v ��?�V��[���>Z��@�A�J�g��T^�
�eKz����Ec�6n)�K��9�MSt��vz�,���+�+o��ҝw��HӨES۵g�'�j��NS���PeA'փg����{tTYt����#��x��x�B�֣]��`��uP��b�}	qG�����6]d��~��<q[� ���X��������S�#���v��WU?ä ��0�=N��8��so�J*���_��6E����"gq5�j�.��ˍi���)�UxR���,:W�kɖi����(���`�Ԋ6�ӯ���/��T�\�%�<�$������5󴉅\���mIZ�����Qm�� 5A��wBO|�_����Cw2Y�T8f��}���z�4d	_�%��rjO�0�vkq>�󭁰٥K��VKj��HO}4�v�z�Ί��G�̢(M�ܠ�����������I.l*)Q�\�V�d���Gc��r\c�XV�7�� Ț�=Y���zm��2(ap	���G"�[�ֹ�p��R��	z�Iy�~��?-]�k(�_���@�KѮj3��I�Uc6�I>�X��S��-�M.k5Im%�I�\��]��D���[�ϓH|m^�'�E����laj4�9�v�M�{E��t��G����7��dr�.z�ۅl�u�jE��+jD��;�6Uhׁ>#�Ki%�<U�X�׷���+��0�5 �s|���dG�q�tP���_dCm�4R�v���BަD�^'{�	"E�>�����0�_��'�~��k��׊w��B�w}A��מk[@�c36�:��
�{$�i.��3ɤ�Nks@H~{Y�|39�x�Z��\z����1���OQ���B�a�Ύ\�6�8,�ԗ�ة{��e��֥�;�7�v�������"G�R��������Ԫ��[r=,�����h�*�u:f���&3��T����ӎ9z�>�xmy.�Cmv����=�e��TS+Vzk`\8�
�C_���D���{�� ���yIb$H�1i��i�g�W$� �����I۹x�@<����.�>�����qNм���a����D��'�3]��h����E3܆��݅�0ް1�[2�X�v:٦��i�	���S�z��vj"�pZ)�8pA-΀
-���q���O.�>��^����#�$(��{���d���T.ػd�%�M��kn��lcU'A}�^�C�d�>O��Z��W�j�Gl��ِ��r1��c�A�������Q�X���,%�ى�ԛ���� ���&��c��_��u��2/�}��a�t0�E��U��Ȱ7;�?�j�[�P��0R���ug��5���N�o��N	A�Hæ�J�)Aȷ�*ν3��Ͼ0�Ve�d��$��EY~!�<�����?-s��Xx�^-#����?i� �|LQUsI�d�")k)�gV�?̰?�ۄ�YN�sfv�Rd{�e���*u��nf�s��%au��蠲�ӻ�=��&=�����M�d���Ô�c"�W7i(K�<�F#�ζ�?/���m��Jt��I�����W�a��ּ �;2�0�F^}�-,v���uKecBW�G��9��5�����s�7���^	���p�	*������#��F[��ê'�(6aSm�0��.�>����z;}R�mw�,�%դ}l������B7�:�̳�2E���u������i��U]}J���2�Y�+SB�!5�H'b�#�P��J��{Z����!����M��cw|���.\����꘬ܾ��od�3L`�<��w�$d����lN��Gm����ь���7*����[��7Z?Ag��"�T�bc;�����?�8� ���"Q6H�ק~��)&y��(�Tm~�<msJl��k`�H��))�8յpK;A��E���w�]{��\N�p~�n?]0�k!;�N[ß��=җ�S���1��{ьU�R�gK	R�����K!oO�Uo'��	;�Wk���u���0L�զ��y�&��1XK����=���C[�u׾�W{P�C_(m�X����{n�H��QA�nu̳��:����=��D�~t��@�c�u������v�/�Vm��&:�3�X�V3Q翤����s��8Y�ޜI٬�s.���uZ?�#^!����PZ� O�l1j����b�	�Q�G�GPpWq�����������"�Π^y(��pDUF<�=%����(���0���{e^0=�6{�C(|� k�KV�I��-�`�������[UHP����]�e�U_�/D �Mr�� ����	�E/�ņL���G�1#���ݍs�+_ȼ�y��sr�@��+f���Oxc?��`y�v܃H)���?#Rں���i����E��,��d����[C(����V�� �-%<��U�F�ȼ�֨��|R�Yv �s���"G|�_v�`��t�5�\f��ɝO���|C)��*�'S�}�P1�w��MZ=g4�,<��\�?�a��Wp�^�i����`��rC�yݵ�XlxVHYEB    fa00     5d0~k�25�0���I����H{�dy:΅mUaX�	�V���W��FrH�)���&6�ǫ1�% _B*��N�{���
Ò�T㨌�*W_pS�2䡀-����^K)z
��^�_J��Ȟ]T��@��e��Ё^��_�nftEyNu�ު�Y�����ݷD_pg�y�;3��?��~)�Ԣ������������eN۪�+�;�o��2b�i0�l��4j't�2+\�����a��H@t����D��6�8a+|��/z�/u%��;s
�IC��T)����IT�����2�o#�Y����1,��2S��Qa�5�KrB˧Q!��T�)0�7T�~8�gG�y���&����ܴ4��󧅋�&�g�=C��]K[߀0n��}�ms8��(���T���&��ʱqH餀�l$�%����,����;d��AF^~�^d�m���E�P��+/�L�*�W��!"rꥐ�����9�A~x8<�
���g[!qID:�6����8k��Jn&/i^K.�d�U��j+1h��_в1^��w09�w�i+䠁�7c,Q��~�Fb�x�@��I�5�;0�����	S�M�C�\�� r�U�*r�� ��uP��C̋4�Fl�]��,ѱ�i��wW��fl�i3�W���/�#N�s,��84I+J;�57Dg���:9=���,� i)�Oi�	����N����)��0��Dϰ?ɿ[�_6�^*ZL:�:���:sR
~�]����C�f:[j�N\��V��e�����M�ЕY��q��zX{Eǉ��(Fmٵmgf#s�9���p�^������\_a6��C��1�����Q#V���h��7ܠ�E�� �ϰb���yn��%y�y��Z���O9���4�w)ţnzP>}H!w:@Y;����~*l�T��'�8`���*�
��/�g��*kQ� �UK����"��v��+�<�^����/K
����#�����=m�:����a�E%��v}�S,`�>�bd��~�W��\�W;$��{M��L�R�bd���a8?�<��V���7��_q|i%tnd��<�;Y��kxr�5�KN��\�q���J�W��<V��j@�No�t��Jn�h�]�G�P��E-C��u.`W���Y��^����!8�+��F`����Q�7Dip|P������G��]�)�%�P6�����]n
���y�x򉩈�D=>{���&jB͗�B��<����_r���O��[������۴�Ǥ`*�O�J��b봶	$ڶ�&�ߨI��T.Dp�� R�u=�����B���Sh�X6�����\+��8�����x@E����獧��<��إ�n�~EO#p��N�b���\���ojjן��;dڄ�S��Q�jtN����-�$@PyP>�%��k��l@�s0�9t��YV�XlxVHYEB    fa00     640�0���N��"�
�~#�m��lt'��//[ ��9�u�����@�ifGCT����;��5wP���]�N���$���Z��*l�=�����XM䙣�ʾy�;��jXz�<�=u�b0��w��������D�6j�3�Aܳ��M9t^ڇ_h�U;gg��w�"/F���L��mV����U>�'ʯ��#��H{KD0���v��f���h�͵c�rA0|�Ԩ��%�����q�/I����T�{\��kFJ��FLzJ^��t䤍_�i�"!�]�=6l��=�:ɥ�Q����[ӑ9��8|}k�#b�9����I<]E���|F)��Zg�1��y��6�藛�u@Ͱ)�TR�	����mm12����_���f9|�`��m�;)��.�Q�fف�y�8��>$6]��"Dė��AjfrI�`c{]�}Ē)���X�W%�v��i�uM\G�<���Z�/7 �w�v�-ަ��� ��3��ڟ��'ï��a�����A�lF��a/�X�Ψ8�C1bAV��R����9�ɑ�_gg��q���S�ăb��ᡸ&�����d���HT����%�Oa���I���t�p�}_�,Y���Eg�����1���A4�'�/u�#Ӛ3�y8rN���\2�x!~K��\��]{P�>���!�9f�H�Dm�ǃ��u�`/��/�fS>�Uɫ�.�f�����o��[O�V���d�K�+�����p�/�L0���#��*>gt�m�G��He�f~�V�� ��R_��}�"�'Y� �OP��bB�A�O�T��� ER�'d
M��N���>�;��X�j��ٗ>~zZw/�e �V`�c�AUg�`�|}��F���\�%Ԟ&�}+�ґ C͟�"Os��hό ���nV�zLu����`Ro�z�S��D��ল���.p�-�x�Sq�,��,���y'�
)�-�i@vtѺN�Hx�]�����2��v�{�f,�$����C�v�y]����c��W�Ӟ�O�g7/�4(a��?E�Vp��I�1�)xЎ�C�O��}����L?�ƴ!�!��S]O82��fMq�C8��N���5��=|��:\� }V������1n�a4�Z�{��Å��v3�	i���������֥%�,�J;?��cn�E��F"b�Z�v�n(O�Q��o�_��$�l��s�_�B5Oם��/�؞Q����F��_�d־(��c�\�h�e`Xs��*�Z\���8H�J�P鵉ˬ ���>����D�>�Xۑ����k��C�>?��`Br�\ҟ}���|LNlM4��3�T�:��@��O>��bn�!q!��n��e���) ����~ppZ�0�����gi���8�����e5���ٌt:�4I?��θ$�M�s"���WB
�tʑ4�]¢W7����mSO4�3�,g� ܋��Z�@Y�55#�.�� ��W��.$���~g��حs�����h1�e���R�����f=�kˁ��t�wI�3�Q�c@�i�m��!�ذ�?�Y�l���c6�~z:��2R��m�0�V�i�j���a�$�C��AY��XXlxVHYEB    fa00     5c0o}�11u-��R��7�C��m��19Oꐅ,�n��%��;u��	�M~}�H*��^�B�5��'4�j��:�fF��u����^{��r�r��xֲ ��œ!�ZI��N5�D���b�l�)�==s�G'���p3��e�9�g�CIEB��~\�rul`��<�a��Ԓ�YI'���/���_��u����<޵�E}#��`ue7��7\�ٹ���1����؜@�q8>��^���Np?{)�P\OU�葲�|\���g��AIfʡ�6��"��2��ZH�\gN&�X�Sԍ=�ۂ�P���N���iY;����"���f��t(�aVb�e�{�ǒ����7�fA�%���a��3�G���;r6R�Z�6?Y٦�n���1�g�o4��?��PB���:4PR�k���P�>w4r7�5���0=����(~���A�K�W�@���M]�����B$�����o�>�3��?�w��� E�C��.S��4�g�?4�ң/B���>��}��P��>���r�r��M��� ��v��� ���;,��4���^�:�'�[�R2z��p~��+(�V�I+���W���,8f)��x_�ϫ����� �ݽAaԱH(P��w�.��.�L��i�t4�J��jj�,�u����9�w3��g�$��F����קFs"�����-� �6 ���ҫ�?wejm��~���HV1�C�B���'n15O��H#[ZЄ�`��<R�k{�`�z���BA:e~� ]���ܹ�`�Y}ܧ�"Pc�_v�b�&_������{UY�S�9�dp@�ݱ��5�UL��ʯ�oSJ>Iz"���)�n�0�@������Ζ��'Z��>T�3�ƫ�,�)`��9���~nh��]�,}@^����I��3[�B�XeoAF23���$%�0
��0s�n��[�!�����%��fX2�ŦػH�i�ė�P�Q�
P���� � z;͢�r����!�h�/����}zd�����^XJ6'�]����xI�W�wg�n�s�aĕ��fb�)P��ᛤ��L��jڗ�d�E;<j�G���mkQ(�U���+9 7��@I�W.Rp]s��B�s>�qLe�#*q=��$ ��TU�x��q�ih�p���~�Q�P%05��pK��XO�J3�%D�)��4� Kv�-����V�DL�?nyX�4���Gq��4�͠�X䀉b��m�gX�KPB��Qп�#Q�E�\D��[�)D *����QB��(+�Uj���F~�ȼ��6w9�P�i6 ��+��.�9�4�=3\z=�x\����7��r .y��n�d�_��M?
2.2����X}
JHJ�7�e��{V��K�����֦�H� W�K�l{|"}h���o[4J(V�n؉#M_�/�O3�|��Vx±L�qy]YL�+�z�(�y�DXlxVHYEB    d347     a90v)V7�v�db�]�����e ��7Y����`�j}�t�o-*+��i<���@�t�v6K�3U&���$�B��Q�@�y�9J�pݭ��w&�i��ɋ�S2��z\N!����4��K��d�9�x �s'�1sͧow�`�1��S̼?͎���ƻ��@\�������ҡ�����rVB3gP����=k����+x��2��C�kpH�i�NA%k�5��_���IGB�Yz}�Iv�0D�t�5��͟���4�,��-|p��y�h����!����D�VEV�`�/�k��%3s�T/	��I"G�N��2�'T�cš�|,���0����%�������UAo�3�!R�	QP�z��™<r��k�T��!����|�� P ���7U>b���ͅc;�>qw�t��!�_|H��
f�e��%�Yrg�����s�F��c���K[mPn+\�\MC]��'[��C%��ڍ�
0�U�E�üWt���
�.G:��a��Vd�����ֻ�,6�����#q��JH�����"#Fmg��o�*��q��
�rq�\(^@�� �NK���Z�!BɫK|9��e{�h�25U�L5Rh�h"����Q��m�Vż�5�H$荏��( r��\��iY\�VuY!��0�"��e'�-�1��g��.��/�qj'��`q�(e��G	�q��E�����V�����&��?H�)�A	����p��/��]��􍐉Z1t�HU���p3�3ܡ�}[�'����Y3O�A{<�S��%�^?�e�]�������\���`B3�ˆ��r9rk,+ɀϕU�"@�-���h�&	�\��4�����Tϯ�%	1���w�+���A a�E�C-�Bh	�ɤe_�u5���h� J�C�tD����qT�yg��7�&b�����4�s�bFK�7]�=��)z���Z�8�� �A��=��Gyy��[:��B[�
�"�o�4���l�{�#�?���ܤ����m7��������������U/���/Ks��c�Y������ ���U$D��ӕ% ���F0��v� ���s"���R]�ՠ3	k޳�B�t��.yy6���qg��J3+�%2dd��HF q����4<��Q��`�����E��������*��H��%9�K���ht��YJ��82x�I}Pp|�%p�PX.��� _dqX�J�QI؇��#zbۻ �͵�HEj�[��;K! Yw�tQ�|Zs+��+9�|�u����C+�pՐ�Y?�Ɓ�f+��N���.j��a�`}W��M�N<!���m߀�#}S��F�ܶ�1˅������g��˼Ѻ%�fQ��Y{>нn�Ũ�{����]uvV!$4t��++�Iڀd�0�!� �I�i���[�u��Q�]��%�u7�_u΍��L��L=$e�%Ԉ�I>�3UE�5�����<:�C�Ֆ܎O.Wc�\R���S�j�9
�rvP��/��W� � ��4�z"l']�t����Gɀ��i����4�"N��L��E�2�߰�z�kl�`��d�j1o��V����Wnx̺�O�멉���]�{L8��w잋�q2#��ϣ��J�s]���J����m��]�S�S���M���<�!�o�r
%���w��.	)��O�P�pǞ6��Y�g���b�X99���޿���f�ҮEJ*�?�/"���+����ðG��όB\TƸ�����E�W���=�x�U҆$�a�l����^�\q�굨~QyA��,M\4�8D�6g��אH����n+v�����޻@��DΦ�HU>�\@K`f��Y�Z����qD���!�@�\�rȺ�ܓ��/M)�1�ꚻ��g��? ����X$x�������"���Ph<�9$j{-�Q����o��(�}��_I��&��i��Ϻѐ�ר!�:�gAb�m�EJҘ����������tё%�?=��̮B�DC
���H�78�p��S�ݾ$ �H�g�U;نMn�<���Ǹ�$���_�-�']*%�Z-?2��]�eFwH��o����0�T��AT�#Z�f��������o����S`9���U�e�m:ѹ�i%ad
�3I�`3o��"�����u�-�v�bm��o�D�C�S�~�8�5�_���w�
T�W�����e(�x�$�lNߒ�4qg	C���Xד�7��g+��qݟe�,~�ߟ\M��>��b$���[H�;Y����O42����z_�zC-��G�V�á��9���J�Fj��S���p�k&��mc� C��rc�"���E{=�t�9�"b3���'Mf��~)&C�|db�$��.��F�6�f��ia�s���[��+��(ĹE�6�-����$�?���T��$���l�� !�������aR�Y���i�gu�����AnŊ���gP�ɽ�}���>uݸ�gs�$��c5�-ۡ0�EqoyĶc��T�i��QC'���#�t�hxgb oK��L�s{s���YA��ny�ONm	3����@tP\��G5�VM��ם�����C]��b���e�^��G�ё��]�xՂ岝[��5��3�3���{�����n�q��B����&O���?��y��_�ێ���O��	@v���