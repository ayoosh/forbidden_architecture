XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���vM⸠n��%�>�yp{h
�s*c��/YGe��GS}4����Ԡ��eF�*�C<6o46Z��PEn=M���%G���t*�Y�� ּ���ݞ��V~~��<�0�nA���̾�tT��2ٽTx���Ȁ���'����<���a�+Fnj���܎��_�y2 %�E=��r��̤I�����fb��9���x�R��X��"H�ƛ��w:�sHà
l���.:�@���z���c�n�9�\
��Bie0z~�Ϳ�3B4�f��"� �\�in�ڱ%��yOl	�k�5,���:�h��M/ڑ`ڱ0�Ϧ0��"в��M#5��`����
�u�9�2,G���H�-�Ke|ʦw��Q��B��kR���Mu5��W��3a���-:�a���r�B�+�$���|%c1�.��{J�V٘x8ů�8�p6{�Bf�Hہ��	��(@���L�⪱�'�o�,��
�c&���3�;R��*9g&{�$��HEV>������	�p�&Cz?��`��c��5��ߧ����"�AtI+�;�+�j���Ʌ�I���~n�ޢ��˓e��_S�n/=��Ύ�#�-4#��/��sb���	A��L�t����p��!�H�o�`��kZ���w�b�t�{��;!��ǌ��*���UY�C=|��^�X��H��6j*�ȟ��Y��G�^���&�.�ad���ۥ��)Z=�JG��}^b���ϸ��ws�XlxVHYEB    fa00    1fd0�l�F��K�ZV.
�C�:���q�щ^����p��|��w^��x��8�83����Ǳ� “����h0������/_�73���Jȉ����9�ׅ�F�B0�(��Wk�\��&>��BL��Ox��^�(�&�A}�$2��@�-֌c�=�lq�e�W�"<  �(fG+�k��D���]��گ �;T=_�-��!$��i�ig��:������̚+��-��lm�h}��%EK�yS�s�c,*_�Ds�(����`u0�e�4|-���^����]��C.�;	{���	��7LV��s����#$�c�E�F��s���#��{��!��:AA�|�i��}��"#?��!�)���,Mx #��L�1���ow��t�<�E+��R����KK�<�d'�g�+�^]�e|Oڛ��[5�Ƨ��T�F䞷�}����Ef��`�Kl#��?�����/ǣ���iX�K7�����H+wE$��b�C�V���t
 J�o�3��A�[���yY��[�qǪ����Iű��q����.��v�A�W$:��g����l\��N�w�
{�Z@O0�iYф	�%o��#o�1`���9k��e�9o%%�I��)v.�6b)E�<*�v�+��PXW_@L�)T�lF�����E����%���C)��������>` ��'Ȩ���`!X�9-��X��&%;���iZvU�$�-.��Р��=*io���M�;��b�􏸱� t����iYL?�w�O���"�җk^lQr~�`�.�.Ԝ��A��1}/`�XL^��e�C���M�c��S���u{�A��I>�m&xL��	"`,�*�3�P1��[�Eݼ�ƒ����X ��⼔+E����pLL��]��0����Q���ۼ���c��b�2d�2-��x/�B��r57�4�T��/������/��7��,Rw��
g��-��<S|_�M:��Il	�� ٬�І!�-����ݨ�i�l����*��L���Ɂ�)�IpD���E����˺89��:<�p�`x�d>�V�|\ [X�7L�m���BY9]M]�MJd[?�����-}���X���H���T"C���s�b��]ށ�*;JE��#Z<>l�ĴSޣ�Z�����~їJh�T�}
ߕT�Ϛ�[2�K[�c�xb�4�\Bs�ߖg �R�	�t"� ����JC	��ĩF���ð+�eJCv��	���|�!��C�����tΔy�$�nW�O���Ʀ�Ә(���Y�� �6_��&�@7hN�R82�!"��o����ş�C�my�NI��s̓��ؒ�yQM���3�.?x���#�&
pz0P{��xzA�}��&K�Þ��'*�����bL�-7��/�q�J܇����4na���8����2y�I����rOCbzc|�$��e��R�1d}��T�.�}8�ًH��_�ϊ��
�A�-�+s�+���s^�۸��!� �}!9�	���%��o�x?)�%f�������3!)�Ǌ�^/�\�����ÔO�w�}�yѕ� ��< d�|��F[Pc{��7p8��	Ml̛׶H�`�QC�B\y�g��@K��5o�����qJ��j��<k��g�ߺ��n���e�n)<�xLh�п�d��8��w�Hh �/�������A�ƿDF�F���uף6��Vx�3<r*^O��nyŞ�v�"1B���-�w�e������(v�  ��s�	F`�}o�[ӷ��4���hb���(MA�Ʀ8��@��!��4��	x������I�G���l N��nk���?�Lq֨'[:�6b�����7tX3��u ��Q6đ�����Hk�27�n����+�0��u�����f-<�sX`��l���֯�6W�9���͍�
L�g���������19��O����{�K��{d;��xJ�yD�H��Y�����x	C��@aș����n;Ȏ�h
R����&[NӟFRw�/���D���y�b>����m�o���eqNO�{f�n�cJ����6���-�Z���}0[ד��ok�NJ��`�H�Z��Ҫan�f��&R��^�ϢI�+�`B�M�F;fk��>&�K�,m̄�hZ�w��w��"�a���Ѱ���P[�PSǨ�d�٩Ók��{s��	3��BB�־��hM�OQ�D�����-���vw������6� }1�%޷�F��ʺ�+���3.�����O�zJ���}��HМ.�"�G�C��@9��s P_��槴�ʒ5R���ћ��Nh������7����0VoC��(�k��K�A>>h�|�:�gҚ��W��|w��0����A��O�QO��������1�Ӏ�ǳ���x!�?�X�]U�n�J&o�N*��G��9�=zp��C-@��F헶�j:��O!�9�Z�����@�~�}���OYM�o�1�{V�y`�0�r����\�F� 2���S��
y
�3�mܲ?�7�2���o����)1$���Z@֧�Д�@6A��(��Z�4t!��E���}v�����1�q[0o-�>��:¼^�.9aW����_�Z��]f�<.ZZ5����A��+L^�N�'�:�Xc���iۀ�4� �V�)��ES�H��j����r�53QF<�!j�؛?�
W���t`0���q΁[�w��C챐�u�*S��Z�lv%԰��z\Ag��+-iU�/(�%(2Qlb �[(cei!�E���p��q��ܷ����O�9��s\G����|�ā+���aƞ�tN��ޮ��H��氒�alۣ��.��9�Z�\d��b=�zh��e����h���-�*Ɂ����z����n�r6p�F#�8��PQ�����L���c�d��T9�鯦�����o�"B	��y-m������B�d����C��@��=�ƚ�8�>�˛C6�|��ifg�s!�����QϪ��}��	�0Š��]%��A����J�5*tw�8Ğ�P�ď�eh�w��퇎xǫ��$�Y},4���w����2��`d�����(F�	�����A5��)�;�l��&�>Ж���D��n���$�j9Be���>����/*�K���(��Pgw�CŠ�(����<�9p&̞��:}�Ppph:�EW��D؆.��x�G��'X�Bޘ1eI�g_�j�[t������[uqAl�$|���X
�;��Cd�� r.q�$�p��O"��qu�ƸL�aϑ���{�QIK�H�;
.���oo�Xϩ�R���q)"���������T\�;7=m����g�V��1
���|&�a���0w^3k�YWv����J��c�"��J�^��$<��$�k$�GM�ʶs\�������W�;/:��J��8�W��,ǯ*���I��>�/)\ꎏ��0s(�ZݰF8e��q{K�B,�Z�d��<���y���'�Bg�f��LzXvA��Z`��/�� X�,����X�K���
�eOӰ��ۏ<ގ�%~ɧ�� S��ߴ1~`�9?+"=6��~�ܤ~���I<�R���9s���H�ܰ'�����z�!H�}�Dqe�����;� �J��M�cx�S\L���_D�^�#�E+�RU�U �}��(�mf��b��D�k��4�y�':E�tso��_��C���_�T X���A�D�پ.�)��^5A� ����	0\��T�I�M%l�<3�|H�����.�`OC��^ሴG����J�[�i�E�Dz�������Y��K{���v��L�)��@��'0�"�S��V�%V��Pޛ�f�i���1Cfl�!��ƥ��1�o~*���طZ;"�l�f��ױ�U���6���z3���o�38�٥_?�S�PJ���.C�#{�2�bR��9`ĸή�IE�j�ޝ�.]5x2�sqY�����A���RG���ƛ:��feM]�hJ�EJ3e�>H��g�3e���℅�c ���0��|Ù~��5@IV�,
a��ba�B�*�:]=��'�p������\EMX/��P10V<l��UVN�K)K����h���}���ͫ(S��U�ݑѪ�
�nN�;�����5=�x��j^e%Gu5\Nb�n�"�+S�)�]�!���>��(�ќ�vp�W���z1&�րr�̌�m�-^�k������lˢ��哑!��Iz�p2pw�P�*�y��m�����`��/�:�sC�LH}���G�V�E���sۏ{訇�f~?���tag��~��ġ\��e��G����:��zvx�S~4F��P0fv�{�̀['�YF))h,��UQH?���oǆ�3(�[ �1җ҇�V���N�x��z_�B�V���<��:�WR+rE3�
3�h%{��T,U��8�=tH�����a[3����o|�������`��حUD���5(����J��~��8!Jp��x����O@9.��k�
zπ�[��65�Ɓ��� �^�􋸰E�H�=_��)�L�a�G��BZ��c͂�V���[mm�&�)�m7�{{��'��q�Tbe�Gl=���_-T�B�gŚn�6�}+��ը�ȲA?9}�!߈k�r���+f)�Q_�X�@U��H�kD�o��!�.cbK���=��K�!��KJ�3�6C(��z�&��؃��N\�3M�J�<)?�`_$">w��r��ҷ\#�����ɾs� dT�@��Ү��J�F̕ڴ���IQ�L��.�Rv�Yf�d������@|����F�x�b`uBk\"6-�+��0JOR�d�G���*�81��|!�����IM
uRXe�N�3Y'tX��=��,�n �V:cW������-v�v %u��LA:y8v���ȩ�X;Åb2�ד�(��/�*Ğt��l��&�?�o��_Fȋ�#���^�?/!��Ӭul�|&��O�������Iv�.zԐ��B�(��D�V�S�0�҂�JRfOz��|В^��@n�`���6P�ږ��()3U��oF����"�<�2�����e!ռ)��� o.�O;5�7ڗr���ҭ%hD�K�F��-�-tI6l�\Djl��I�ч��GK��ʰZ�[�X� ��Zߙ=7�|V��x���ZE7Ɵ�D(�}|n�{�c��D�R�8S:#��-Lg;ʳ��ПV�修�6����VU�z|s)�˿ή��(��@[����)/[��׆j匍;�B�	UA�U:FP���o�4҇,<rE`�g��fn�V>��l"y��zvZ'�{L8�}P,f�l=YB��v�*����X��dl�k��b����kt�$(*ḿ��\yՐ�c�%�RùEk��_�j�vި�� \�	chA��Ͷ�j5\��כ��G��8�e��$Z�g1�{:-r[(��t'S����R�$�;�P9���ߋ�ưf^M#�D���;kL���8j)+��`�k�SCA���m�A�N9M��Ӡ@�N�KĨ�BӚ���m�\M�_TxTO�ͫx<��w!�{���n���E6���q�/�;���' ��.a� ��#��|dI��̛7=8ET����^�Ū���D+��.�e����[�gri�<�o�H���{R"d��흾��y�&��O�x"kO��ZYKZy͒�k�ZҔ�Z��lv���?�ř�V+��@2*�j=�� ���̩��]���F����e
l���1�c/Q3sM�P䴗���#�߁17���o��@39����'e[5�nzZ���nG`�w_R"�Ͷ����^7qr������k*�h�s9Ε2Y(clc'�:k�Q-�'�1V�J�4�\�>2_�8�J�N�$�fX�q0�:���
�� 5,�=i,Oe��	���F}�5�,�qk��z�v��Y�ؽ���+�7&I�l.-�~ B�>	�*�n���˯x�U���i�YX�lOd�i o����K޶$l�ĸB�b�hכZ!��j����S8�"��(QB{'-&:UVz�6j5�{6��I�"0�N5�z׵q��R�(�Ί�$�y���/�1a�GlU,��.�
3�v�o�
U�m>�JE?	���_�H|%���k�%Y����v	��+� ����؅�:g��[H��As�5�iޔ��lB�[�G��G�@����G�+c� ��b�Rܙ�^�XڹO���P�Da������M����� ������������\(�<�EV��8"�W�j߾��$	��/Z#ܷ������EOم�_MR�.4��\�Ko�)��jc��9Y<�+�S�O���)ؘ#�u�03����m˗3a�M���~�Ac����NOy�����!�)��d���4rKn��omN�H�Rڬ��=�b���T�fl�_��0mҬ���Ь�	�eb�p�t�L�z:�p����j�y}��d�=h�>@ޭ���2�fJ���=�����$�רd����	��`��.�X����%���A��Dq�	�G.~㩵6k��2�	��ʓ䆴MEĝR���2欞�q�Q���3�3U�#j�x���?�\A����F�ܚ�4LE�RZ8n��a&��<��j��$�03��d:(»\-� �e�<f�#т��,S�������η[��Ҵ�R6���*��+�?�Gt�{����8��f:��$L?{��?s�r��yN`��p�N��p~Z�jf"���f���\��<>�ۙ��B����[��}��
�+; J�	Qᾑ���yfE����@�k3NQ�.�?�_��<8`Z�S�QJٽ�|?��������!Mu��_�=��Ʈ�)n����xGe��� n�s�Xg��X���o�`f��HRQ���W�,��K�7�H��B�5�8�Q�8��ҝ����fӾ�>gދ��h�����z�s&��H����,�U����*��i������u�\DV�%d2=�M�hm����(jYʛ�:�y(�Ȧp'U��O���{��i�L��lT��ẇ_�e'�]!$�m��)gh�FNi�SD��+H�{#��
d���mE��A9�������"�<���Za��v�p�xp+�����9U��Cv�i~�=�� ]��o�aj�M����cAi@r"�1:��Q��s�g%N�v݄�����[Ę^+�D4��1a^�<��^��I��*X'�AnM��Ӣ������Âw��{*�eQӾ��*KcT�<�� f��UBC�y�z�2[��@�M�=���d '������(���>��9\����DHdMyۨ��E=#�g������ܫ� ��pQ�L�Fw����׻$�?�[�yR���S����>�Jc�æz�[W�kɤ|"��3Z�ʁ�=��x��o����zH-Ciw� ��4 aekR�Z!NFϳ�/1�r*}�B���:��g�����7�.K�`)4�A1��\�#g���/�����y$Y�z��xPRm���'�ѫ�p\(q�ha?'����cG���G�y8�jACLot��ϵR���W~XF�����8d�[���?��o���퍏{n�-�֫��?�(�b�ڣ�E�=̉~Y(	�	k��;"��7>�ɵE~�(kʣ���!���Ȃ'e���Mof�#� N��i�K
%�V�r�Td�a������r�����8�Vs�d���-f䤰�F6���+D��ja,���#7�2�^B��+p<�q�>��\�)�]xI��p�U��S���(Z2�҅V�����k
�  ��\Y�ۜ�ۡ��9����6?m�̯v�Sy�V��A*���`�
��@G��
jX�	{�>���!<c�vnH�7��d#$��6"O���� �'�sd����L�ƶG� �e�S��B�x�2�@�M@|������흫���c�������|(�]���)ffK5N�� 2�Cx��u�\	KFA��#��
���d�TQ��.�����n�<7��[���JX�j�������]bŃ�u��Չ�W��b֨�n@��3�0�W�Sun�p3O��=� Έظ�i�XlxVHYEB    fa00    1340s:������}�Z(!��s�� ��zMN�kQo��F�V7�}�/l�5uNM��A�˼�K�x��e�I����/�{��� ��$݈5�h����A?E�~���V�͖nh�dR��j,�4}pm�mF���y"O��qoJ�E/	}����Y����Ly��M���*�h&saV^Uk^�%Mᜨ6294''/bq�кmyt���VĆ��9�)�A�g�}[�iD8Fp:� 搰qV���ݱ9+�0&y�z%�k����>��'UF�3�uμ��ۣ��%�%�_}\��hI]"8Vt�.�#��:Q�g�~k��c䯅Aܲ�>����S���<��K<�C��O�	�?�ਫ਼OG�qj�p$��vȝE5����<c�)���\Ong�6�4ٗi�I��x%o?�ߤ�w�F���,���?f�(�(Z�j�d�ጙ&J���g�즿�o�d�d}��,^8J��\�
M�J~q ;��J���;v�y
�����PDu�O�ֈ,>�^�Z��4� B��~ҡS%&G�ԫ����K(1��6G?6Xzgf��f'e<����.�t�� �p�,P������db�(r	7���!C�8C(,����wӏCd~:�G��{$ˉ��)�󣘆�����P�aɢN�e壑�ʉ�|`�;�� ��=�4�l�$$��<�����ۜ�����_�	:`�Z�����FZ���ƙtK+��(��č�ꮢ��1�S8�Ip7��u�����+�'Xb_��1��p*?�w�auB��e����,ET����e���z��Ѿ��g!�{LѧR�&�柗SN�mX���5@F -���}��]��=����#YDz�)��ʃO��;��$�`�9��1d�Ut
D�`��$����u��g��y/U�l���Q��������Ғ��\+&�\�4�Rl�i8%��G���e��]�:�m��-�;�
y\,��J�y�
�	p��oP�a#�	^������U�7�q��ތ�ۥ�N��!�/<�W��,�<�l�{õ�_(̓��I�]c�}��2^�l<�F�7���mdHo'x��~r�����s��x4�V��WP-�Ez�h�[���Q��eVIr��z���Ā�s��,��j�05����L�fJ�+J˗iM�P��:]̽_^�@�&�}XZ$���Η�;Y9t[?Cb������l[T�N���Ɩ���������k<�MK5�\��\��K�(�l$�e�C�3��1m�_�����\��S'{��4�}8SK���M��Jp��8�ʣNz3�(��5�o��e����ޓ9
�ܭ{Ne�j�]w�|��V����)B�Ji�5ܻ����k��sĨ�u��@�+ �)�������v���"��ōu����Ճ�8>�H�OaTf�vӳ�]�{�)��x�xGޑj� j��{���c���}b�"�q���� Yr3N�;0�1��s���e��j�b�I3�2�b.l��ʩ�W�oj1���� (R���V�l蘵t�p�3���q�&�w������0� yCe[r�^��BH5��D�� k]���8=�*jY����9�]N�z�:s�N��v���7�e�h������+�S���m�����	+���f#�mp�y��]׈�e㠪��ry�7�W+���n�cSO���	���&`���F��8�� Ņ�I� ���t��Yu݌d�UN��D�m{���>�}���k�Mp��;�t[�PC�wx��s�8m���ݪ\Ez,T�&��`���
��5C7���P�9#�`�~��$�ۍ}g=��u�y�fG.��O
ߛ�춻�SUh�ټ���'��t֪��;t����D螌E8�Yۦ���w�QAM"��q�/m]�q1��LO)h�PE���Ug�c�g)��C����e�#�V��Ϻ���D������9(�B
]��M$�Kk��Vtm�a��:1��F�j�#B���ґ�5w2:�"��C!ߙA��)��(��}��̕���s��㓟`��N���1��-� m�M��&��(��m�ϥ�$������V8P$�H(�ם	�2�f2Ӏ���At�=ʂ�\ u�`AGh��՚ס�h�[������a���a1%���k8�#�m�:�9w��Ѭ0H�����Hs���i�&?��5k�;i�삃�i��yUmLV��6��S[�e����cO�/�ҵ��q������*8&Vtű�N�@	��f:���um�Yr/ s�7�V"4�= ��q������Sqq�w��hnw�!`q��+` P2����z|�1Q `X.�9��#���Oo�(.T1mb��Ќ\4���}�����Q3�%��ě���W���2
���L�,B�`��}^,$��ˑ�k!<-<972bse	�⇕G�W�C��av�?DP{����IC����SWo_�ׇN�1E��(Uŗ+=C!E��eA=�r�Gr�k�%L�ߗ�ǚ6�̶c  ꩪ���d~V��_ߝT��]�3��o?�ͣhD;M`��57Y^wns5=Y��S7x�쎨Ӧ-˜��ڳ�Y���x\P�jWi'"�LD�8{�8��~�����%�?�Yj(i��ޞ�2��	�>���W�d���A��Қ�����&H-�b�(j�?���$���M��;)�ΰ?·R�[9"-Ů��/�̲<t!y�������ޞ�:6Q��z8tI��LMY$:1��_�ZJ�UA��V��d��c�Pwh����|M["1�I��� ���.�}�&���>�pLj����) ω���Z���\�ab�8?P����a}m��>Ѧl�,���m]�$�ȳ���B�6"%Y�C�H9W%E;bU)^x�Q��ޢ��V�R?��q�7�꾃��b˽FٙV�Vt�.7��oؾ���6�5����p:����O�],��&���W�m��u�i<LG� �4�I����Y�L
��i}��]�j0-� Pλ�w �/V��b|fi#�Fbu��P�uN9M��^�j �}�а�E��rW�	(g�;�u����`��ģ]ȉ��O�gyX�=pS]�X�Y�r���M<{W����K݉��.��[���d5�x���ݹ�4�Q}�.<��f(���(|j�a-P2$�,�����C�8y��� zZm���a��<�T�?�g٩D�s���J����.�d��Z��(��ېb2�r����,O��m~3%s�<no�H�.��M}�G�0�WԠ_�'lm�L�#��Pa��gN�ǐo�K�2���ǧ3����}4ϯ�-S���x�~���yw����w`$�q1�'�O��b�6|S�U�4�������;��_1�����.r����֊���n0�mVP�8�4ȌD��,��O`ʇ��#��i�v�p㪉�s9n��YD�����Y��{x��X�����rK�wHL����t�������B!��/� T+|C�&�!�(�%� b�]���L�v�H��
��o^uI��=Rڣ0�8�e��d��4s�\XIh臉aqM�����?��q�a�w`� �6�m}0��@���J�����:�?md@���(.�]f6S��͍��'r �g�8f�WVm&H��f���� \·��X�<��-����\cC��U�8��	���]7���ژ|�#.�ucj���
e7���(Q:b3�M��E��$9��g���H-K��U.}어��P>q����%$+�����yQՉ�>S\�#cx�uk՞���۸	���ܮD�g�����c���&P�s���.i���L�2�A?��)�	����B!��231������.c���ϔU��}��ay*y�F�ȅ�0��KL4�z�sQԓ"�L�Z [!��5ޛ�p�+غ�K��>���Z�D�x�z�7�B	D�6X��1T�NI����J]@��$JL�:J���ݸ6����m�hs�E��s�@60"]t������Q���CDw�;=e
�*�����+��1w�$2N&DW����ק�m�6>�a��)A�������I�6r�f����n�RJ�l�:�K���L�j/X��>��C4&���_�i���+,��Z�z	��J=C:�y�s�:J2-[ur6�:	��ҧ��۫�۾�� A�/��x�/g{����v~��o4����c�V�'.`�%�w��b�}�'Ɏ��O�2�pNF�6�l���:�h���e�#b���*��W�b�ɿ�g=kY�~6�%z���['�����nFd1d��7 
��3lFX��k�[���.�65���=�l+��}��J԰����?!�?�Z��Q��T&���A��2�2kP�s�6j���rE઼�f$�cD��8��E��'W���6J�1Fi�= ��J�m�S���<���7:yM���o�$�R��_L.��!��i��#A�\&R�����[8�����g�`/|���v�i�m�+��^��G�Ӱ͌�)�#��{�ރ����[SXors~%O\���]3m�.������ʼx�����n�8Օpw���ag-��=��9��d�_���n.�֧�x�8O�IҀ��^�V"1}`����G�C?^��N����x��	X�6�\��K��Z��k=������F��U���}��!�����w��s� �N�JyZS?[C����P�Xӗ򑅾Yv��58=��a���DV�}������J��?�LX�NRG�����<��[� �[q�9�-W8Ub�~��A����F�'������	���:�)�r-K<0��z��b����Ũou°F}XlxVHYEB      e7      a0�:TA����qԡ���K��g&����]�~05ўb�^��{b�D�~Y*��iE�9��n�!�":
������������8z�fL�"vu&3j� Z��o���\PbAI?���`�rbA��"��tA�M5�W�ȿy���/+��,�z1e���]9�)��