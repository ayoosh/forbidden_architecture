XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���d�՜�ם ��c%/����K���A���	rs����!�P}���FB�T�[сvS܆�
�+Y9��d[\����)����,�I���8����ɮ�#�h�4�c��;������1�z_N�(9O\�3w��~ra��3V=ЉLHFOp6�N������G�1g�Ӓ�'>���G�-k	M�a{��e���}C��wت⭘�
5��y�-�ȑ������|ć�<�����y����S\��	�9��xg�c�+�Wry�W	�"<�����ɪ �@��I�T�á�	������;�F�}���D4��e�?W��*�
�L����5y�������?�n�XK.��
���>��6̡��s��sH"�d1�Ado������(>&^�<���4�+�d�%�����S�$|�N$}9ֵ��Q��+�h����1�a�b�ɇJc����H'�����z�������
.�/60d���_%��p�#�U�;�+����umIQ��	iI�_x�o���-�j�h��6�4�j�.��=�7�g�����@ږ����1��'�����*�/�3�c�W�rϴ�T���rk�N�r�h�Ъ4�Tsvہ�tPfl��@����0!�ql���)^W���u�:�p"`�e�ՙx[֟��z�)���z��m������JK@�L�q���L/��M����R9~Ed!J��USq�1@~��pKɳ�g�A��#2V���#�A�Kf�#b:	o9pj�XlxVHYEB    1427     840��Ή���Cˡ:�����
�~jVL��H��薔ģ4�`[9�a�3�SÜ�Y�����9��X�0Wg�1�šSp�ލ-�Y�V�X'o�*���Vv N����P�u�=�;ݠ'�f2D���^3Dc`MY��6�ύN����'�忦BV�@�QK����8]h���XkM�b�sj�Qx{�٬	� ���������(jya��<wP �"���j��B�z׮�ju�xl[��ҢT�=�Z��p����� �6+��i��l���v�8�hRph�Hz� ��Ď
���k��,��u^PK�۳� �:ģ�D\��UAA�G�?�>ڨ�q�P`T�	8}6����O�w��K?��Mg'5��}�<�$B�\(�I��1ẅ́�]*�A�"'��DE I@�t�:�!u0-e��jM!�9��6-q]-���4<i[s�T�vΧ�G�Ϡ#�Ҭa��$�"x���f�׍�+���~]�+���9Oh��t����=1���T���Δ�Vx����p��WUp���Z�Ŕ�k� �9
VS����n����o����Bl�G|q��i�g�E��K͔8�������Ա������|�!�c�� ,ϟQ���2�ZtUT�q�-M�,�;<���v0�Qmw��k�Sԅs��h³s����J���L��iB,%�cٯ�_��Qׯ}�(`�&�?�d���}T�N�[COb�ɾ�>a%���S J��z���%��.�����u�N!YL>�_mM�lIsU�̾�i?���!�<X�
��ȿe�[��L��hv����l���4�i�}�-���v*M[YB�v;�Gv���+ȡf0?�ݯ���hE7�Ù��+��|���GNg-�h�=��O�>`.
eܓ�/O��Q.�%g<�hy��J���b����k�H��L�A����V���5��Z��I�~#H��/���^���p��P��f ��F�o��mg+��u���`Tֿ-W����I0,u�R��#N���%Ipa�WB��L�����X<M�gs�k"P�I<��κ O���H�sԎ����nS���d����@˝:�ǖ�����]< �T}���j����/Ȃ�1�B�V�b��e�!U,��DB�D}\�N���BL�k/	X���Uo�BU��W��u(Dk�
rj*k7�8D�1����c5��N�f�0d�}�̘ff�,�#�P|u�;ǳ�RpRUC+;D1��s�1o�K�3�������Z�#̆���s!9�9�U���E���9�7����τ����+ĠR��)?�(KH$WM���8y�����0�;I���ؿ޵��1�yu��S�ɶ�.��DQ3�Y���i��bc��<=����� Y13Q�)�-$��xvA�BȾ%ĄB�4���Y�>����UE�6K&��JLAN����١耋���G��F*�R�Hn�f#��d��#�wK�Z��O�����o`�>?ǰh'EZ"�ŷ9ւL��\�ÉJ�v8�DX��`�%�7;��B�	��AX~�D0E��h��!���ۉ��BF���Y �䛹�~�=����H��
<� ���m}k�3*����������K��������'�Z��G8YG8
 ���9-��T���A7�=����޻��I��<4�Y�U�cs��rZ�<���b�XLA�tG�JZ�"+=�Q[~�D%���I�mH�n�
�-�/�dY(
<^h�E���4���N*	߾���@{̫�J9$h�*�_�[H�9���"#�t�ž�?lN'�˳�HX_@�#�([�׻l7���|�,C��K��H�ڏ%��o�'�`�)����	����.��)RQQ�����1���7�dߛj��� �Z�R_��FC���\oa&K������+#���F��rg4�U�< g�'sj��	Ѣ��l>����}�֩y��?�9 ��0�8կ������`�$�-S�0^+���!�tS<�!,����Ak�Sp���~�g��E�=o�<��!'�2u�0V	����V����Q�`��f�����)�1