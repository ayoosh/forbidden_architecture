XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+)#���-��^})�MBb��$���v���AE5D�j$F=yҷ&�js�΂Z	#MnbB ^��|o��nnZ\+y����}�0%Kµ�QA���:�,��Dn;v�E*0��rB��ż�{�7�����$��ǃ��
d�:��)��-jB`�(-���@ҿ��:��]+�q��P���5���l�2��R�PA�᱒���?&�`��,����G��K X�����h�s����.��K>���1~Sg�ձ�~�8�fO?�]�BЯ�۾�;zΪP��nHH�� �Z�;���KY��jQE��(��<��	�ݞ�ii��=��]R� DY�A�� Q��K���g7ˤ�T�SzL3���`j3t��S���1[�6=�)�c�n�}0uW$*���Q��.������˿dKs�R�	�G$�;K�M>3r��\z)���/�@@�P�b��R1IA��f��������Un��f`΢{�MB�̢U����ɳ+��B_B�_���]��ReݭI�R*�����Lo!D�S�]!��
�c[r��&�5<y_n��]�Y_G��&C��Pi����c��<ʿ-#�x�7[���`O���4�lKn �r6>�|<�ʇ�a��pU0�N�<Y߽�%��7	�h��� ���F�P�JC�CC��-t�>3(���wh퀈�/�����m0�Z�Yv�a\w`V\�*�k����#���d�A�/�+Ќ;����Ĭ]�J�l����1���6 8d��XlxVHYEB    fa00    1790�è�"�	
�� &tZu�mR�������?)&����ȁ�汣
���ͩ#̷{A��ƾ� g9q`�XЬ멘�-�V��Ȫ���h�ٓ�����dӪ��J$���CE�Ri�k�I�&�)S���d�bwX�(*�&+ӁA��_��ZY�A��R�����(x�g˴\�KF\b���)f�E���+}���@^����"w<o�=p9c�:̭k����Ľ!�����zt�s&u�΅��"/���C����%�0�!C���j�or)�p ���$ .u(�ڥ6e���_�a4�7�i
̨l����Dl��g.������y]�9�i�f��s�:�ҫ�������g�<B8sK%y��2Ŀ�/�~vs�<��Jy�"z�x�����Y����������!�Gz��,�Ԕ�F�!\���ߊ.���u�VQ��<���GDV6BX�zL�9qۖ^N����.+Ό���m?�׽�3��4�񡂡�Qg���c��|�|��y�Q67��{����flF)`����t"v;��D5p:��<vM�°E��k�]�=������K�C,��8~ĠA��c�$6	�l��(=����\q�l�y�Kޚ���ңiG�u�tQT�n�n����X
e������Q�oQ���څ�_�+V6�R�6;�����U�����G�t�,���)��E�3Br�2@C���]H�F�����;d����]�\<�֌fx̃yX2l�32�����q�ͷ7C���Yan�(fC�*�������BV��P^�D���0!s�G�� �1�-�ysB��f�*�</H��_�����0[G�+�u�_T�e84-��7I��;w<��V�N��ǖ:=��� ���Y����)Z.. ��UZ���)�(�̃��^�^ 9�9WN������0�TP}̋�Bq"r(�A��h�#_�U�� ��|ֈ�!�4iS��H�)~��s6Y��gK��2���������T=���-X.63E�e�L�<&5��wc9�ӆ��̵^����kS'�2I ]͜�Ȯ�)�/ʩY�߮k�^��*+�b4SlsX���Vw�)�ɮ�k�kے���^��>"xx�i��^ �`�!7i��m�s`�Aט�h-�
gH �.�2���AP�Ed-�ʂ8�/�	��Y`	�hPC�O���S�Z��/�Q�V���z�� '����j	.�>v)�Nr!��˺U�%�ݛ��Z���"5��s�~�ay	0`Ξ�,�e����
��Km|�RAk��v�� �S= �eC8�X��?6{z��n�7�� m$'���I�?�[� q�c��K���T��S�Ӭd�X�˄��eG��-v�U<�\m����?_�X�Zcq17�S[�5���?��5���%�Z��9��@�	^���X��c�ɠ�ϣ����R��ޣ�H�4��'�1*RZW��34&�[�k�x4�.5� ���Tb�:EדBE��|0Myɬ�t'͉�	�����I����_������'��)/��Eo�w�5�B٩��ߔ�P�����h)5���I#<�S��-{���ʅ�g	/d�R]��YC4��Χ/lx�e���yi�x����ze]�wە��>@�G�����Z�_����m�v%��L��e�ޑ����ҙlG@����gT�mnx�F��.\i�n��/�i�ba��P"V�h	q�KYG��wx���K!��)��n,-��s��w�x & Ih�s
��*V8G�T%a�B���8���G����-h��^7ݓ��)��� �^
��+�l�!m�S�����[S},(����O��e0כ�v���0d�f�z�O/���2�sx��R�������g�WvMo�r	�n�D���L��\8V��$0\!�1����)��8�yK��$�1�;���r�J�r���.x�
����%�}� �{��f���QYI=۳�D� [aR[xI�{[�m+����3@
�m=ϟ�/֊��팭��x�j���
���(�[�Q��UZ@Q<?I%��!=�uR�`&r�9�rf� �U��jwYx�ë�te����%����x�'OXj�|�i1ta�|�<UJW��;�Wp.����n�KQ �����<\�vj���J��)<� ��Ói�5}����#�Wv��a�1���eN�<������O{�G�9
����n N���f7�,���5Bm�o]kLIb%��x��� ~Z�^󆡭�R��$�}���u��JB�ۓn���X�LEEЀ�E7!�P�Ǝa<[����ц�0�f.���V�}��HK�<�@�����3�Le2S�;nۘ����a4V_���u~�RD�YR�#�5P�s֫���̪�n,��usO/����aBE�j�~�SZ�JZW��� ��}�*��-h�4*m3?��!�h�
\L(z�:9�!߁N���i~bM��Xm�-�'�n�;���"��4���es;ep�K|�`��w�܎��+gQ�z��z�o.H�Q7e� ���}�f�;�R�n���/��n=1�XO��5�?�%L��o)��;�>ׄV��x��}h]�h��w�M�
��ų�y\Z?7�i�?�,=`�i�n�#��O����;�O��a�P�*�Y�^,�|Y�������`&��r=~뜟�n�k{�� �H�'w��_eD����Y�!vݿw�7��T$��2�a�r��=����zqx�(G9�=��b��"B��/��]dx�0D��Le.m�~�&��5��b�J�N��*."��G<g�%=�`� �@��TM)$���b�,C->��n�����#���
 �����iؕ��fF�x���J�^M�5Pc<�����Ú���Rᖗ7����� 煦P���Z��S:ʑ�=/§4��ŉD?VKp����p>��I��K�¼���.��D���U�j��L��l1c���iX�V&8ol�?�}�kd1}8�R}*�,mˮw��!V�k� J;�թ�u̹���$���P6��|S�<�֜<��F��lTϒ�������m�����@����(�Hg�t74��T�A�Gq��5�����t�o7d
�J�ںR?��-���r0 ��WK4�+��cMU~�� x�	�fQ�:~�~M1����إ���U�@����gz��ͥN	�^$ɐ�����Z��6]��e+A|�9R�-����mf����P�;]X%j�\&����U�����M7Є�Ƃv~�M�� L�$�������e�q74����p�i�,�(�� ����/Ђ�� a��c�iԴ4�aG��%v<�n�fy^3QA�͆W�*>kW��3�fE�Y���`@�6v��b]���e�8��+]�i�W]�ڶ��ӎ��d���h�`������VQ��2t �%68���!bk��P�I�`�.y>�}п����qV��mf��O6���t�D��n������P�(�^�yǆ���"����S�G��0�E��ߤiH)'�I���Qb_=��Ko�=_��zx=EuC�S�`|�>���~�)��(�a����r/�L�\�k�.����l��}J'�|B)5���w.g$���j<����S�D��S���\�Ķ`w>Cq\iõ�KT����$�O�P0�BJImx��!B�(�~�6»�aj΃��4��}wcd,U�A#�|�mbmB�˖�c)��������[���#�j��û�n�?cup��jfؚ�c��/=�!+����4]T��q�g=go�4$���	<<]�L\�S`ǙM��e�u����)�Չ��a��xN��Y����Htڱ6'8�|{$B���tW���U|',���wz�p�l���&�d�0����vK�.�(M����{�I��'Ǌ�������@T�Ku=e�o�ٻ����;�ym�ѿ%K�b*;L��C�' [���Jet�۹��	�+� P�1Z�
�*Ӓ���c�B�H.��� ���2(���Ⅾ���`I����϶�V�H�mT�D��A�f	o�->4(��'�����c&Õ�=GO�mҘ�*�m�O�س�"�8�����y�Z�e�6�&Q����l�0˗2��;�E1����f
����8v�bì���I�XG㽊�3�o�(_�LY���w�b�Ae۶ q��W �#3���p3��'G:����^ T�װqj���7��*14l�r�����B�=��讀4v�hֶ�Jb�(�f�Q!����6`�A��Qd�W��� �t�u�[��n>�z%
����U��������4tN��Ԅ�i=e�ӧGJM��\:9��6��o�J��Qn���ѱ��װ���>m���a��zW���a�d+�wwZ�!V%��/�7������&�����2$/ˣp���c�y����f�^��������Z�yŞA�'$|^��jY��M�1�VY2�3�ߑ�(V]�栔W>���m#2�I����w�}浢�"�-b��Zk4[�s�E�@��k�.hE��V�m*i\�.��.�"�)�=���۩��r�s�>�dS5�����_羺�|ϩΟI5���W�s���ea�|��nzg����*)���[=;��e��S�K�5�߳�>r�'���n� t"�:�}圶�O��R}*?�Q�O�����3�%)����;��UbA���g[gyxټ[0o�5P�D��)��Pa<�x��y%%�͏{������sqn\h���_�g��=fg�2���zlo�t���,p�Xa�oHv���UL�J�]�~ITS$R4 ś��E�eq�c�; 8�C/�Β�P�"4��V]���3"����?���t�|E�)wŧ[x��3�O$W�|�_�ƙ5���^T�砩W�s `Mc�����"/l
�x��(��:�r�Q>%��wPDW��Z1Q�h�#6Ř�~�e�B��9nMb�.��[n��j��) ��8�lj��p,��q4���Qf��O=��I�(1I%�&�\�Y�� ��K"FC*CK��b��`���)a�dnZ�ͪp�#8&�7ΐ3���p��-%��ܼʊL㯫a��$��)J�x��vd&�6���'�2X񦲎V	�v qCQǙ���;�����\��ᐹ���c�OvS���!�;�~���Whӵ⡳���tR�#*�@
�E�f�uW���{F��g�}Kl�?aqB��
�s8�W\�pJ������+ެe����H����A�[�)g��H�<�VY��0�Yz��tJcH&�<�L0F�+�wdt��	�O�cs'>��1< Λ��gt��=7�a�֩����z�~{a�C+3�ɻ>F�_3~��Z�7�9MP���LF�Lz�⁑�v����+Ǔ�Z:���v�KAt�PԾ4�#�EV"��
�lIx��f�E�79��_ ��-�r!�d���	�y���Mu���+f"�y�'��,�؟6Bt��p	�=��Z>}5I�~_���)��Oڥ��0����~HF�`?k�ji��l�#zwl���M�m:Iq���D�8�_(��y3�5Q�r�3��cW�[��#�"��S�m�~q)�l~�c�n���b�I}�MvĬ$[� ���%��-��D>�e��pU�u��A�� �#7��vV٘�t�����}lb�15�{��<yB��E�ץ�'i�1�@d�)�_w����I|bᮛ_�m��J/���������$�ђ�Xcߗ�kɥ��I\097�{ŵ41�R:I�T(��-
��v@C�>�vE�s��g��3��<u'v�YA�z���}�RI���j��S�D�yf�|��/�9�3W�)o��"��
4���{�:��g	|�%5R<��� k7�S6l0�$w̦ Df��Qbm�ކ�����Lzda�a��=E���r� �[0�5?"DXlxVHYEB    fa00     5d0I�'{���Hb�{Z���ʀ���LY�á!�u3�9|�y��}���S]�6@C�	�v�_Mgk-g�a��؇�7���KC�L�-tm�x |)ɸ�!/L\�u��x��b��rQ ��Q�!E���ɼ6Kst�D��� �ƫ�cCrevY(%�����!�j>p�nم���Ex�F|I�P��$�xQ��:�M�P���"�}��a_���5�[��>��a��#	��ͽr��	��ӂ�fr�0\/�,�a�L��?n�F�v�ޮx�<�y���cڬ�%�!U��j�3F���m��7k��~�̋M���R���X���V�<�}E����������l��� �k�#�W�U���7U�KJR��mQ�*`�����JT[�S	��\�ص(i.u�������Y��!���ѥD �K�ĽB�-+r O#����P���-̔�'����^�ŨfU�h�/w�#�G�� pmT]�[^�X,��4Ӗ�ɸ�f%��_j��ƥ��10Ioq>t��9R���l�[�������j�Y�V�:J[�	�����
���r���V���l� �lD�ѩ�Y>z ��W9��6�|m%��]ۏ��������X�gh9��e�.�[��uu%�dv��ƭe��+�b}7���"A#O��I9+�Myky�\1d�u��!5�QאK�
0ˆ�8�k|�%�+��B�_?1��M�wVj�5=��Q�Ҷ(ǅl<�pvu���~&�w
m}ׁ|���9�a���o�����{��~+Id�eP~��M#�+jFg~�"d��eё���H��}di���ϰ/��<�t�aS8�CAF\wȡ�"�<��@��7��@�Q�\6��/w�3��U��Y5���)���ן�As�AS����9�5�{�ߧ�`��ӽ]�����*G��F�abE>h��$8���������N�dd�y�D���! ����ą~�sa,�����]�������,��=����~��q~4�m�J�p��(㒧�UY2�FÌ��nU��y0����N�"�l�N"�R;��靹|� g9L�C�.�q2Z�6�C�S���E���C�e��XD<�3jV�,&{�1q�K`]6�P���\��/���_�=:�(m�\����+z ���vkꪂ.:�-x�f��C�ܘ�i�'����i�����s;�N�TS�,���ߊ�k��K���_�w|�����R��s}���j�r�!5�Y��|�'r���g���h4�E&�yC� 2�<�V��d�-@�� Z߸���'�Sᩮo�'iJ7��%c`q�ԋB���61udW��� ~G��2���d�����3|��g���!�"Z���)����p��4i�(iGC�]]��S��(�J;쮡�^FҢ�_�o��MQ+���\�:ة�"+�z�F� ����x�G��[1w��QM�V^_j
��mT����E�7^�Ylˡ�XlxVHYEB    fa00     640bP�GIN���l$@�_vo���^�Lx�|䕐/�#_�����N��@�/�)���hc�f^Y�Co�U�L]:V/#�����j���W^o��е�k���bË'8+�H�H��%�W�M+|PQiBH�!�I���>u4+����	��u�9��֡�@Ꮖ<��f$�Y��&���޽4)�]�f��3�q��oc6��#5��_[����d ��^��U]w\���J_��Y{*
u��	]l��6_�H��K��)�'�L�_��L-�N�$�KNC#q-Y�)2dj�?�@���T�n��t�J�?��!���tRS^c�:�A�S�L�;��]��h�E�@q���F�L��^Ȳ��J�֑/���R?Oqu���:tg���dz-�$��!&���������	_�[/V_Z��U�I��h�'h�<����
P�'u���YE��͟QFj9��=�u��w�W�lz�(roD}/�ټٹ����-^����	�Z��A�/c
�A���1	��%[?�I�[�ڌe��=��d��"�^�S��^�������'�2g~;��s���6��_r�CY����8K��!�����fm��V�T(ӑ.�J?_�ǭ���I��6]�n��qF�	�{5(㱘P�^��V@��=%D�!G=���^�yN1��u���<s���+�f�=
�AZ��ho�{b1x�v�@�wQ�s��nG���;-�5�v@�K0���H�����?R�F.�cT�`��J_���̋�B�('�Yo9*�eF%e��9D�t3�,��C�E�N�J\��aY���g��֜���H(�F�8�2Чh��M#���~Iۙ,O2�����n��|18�TZ�i:m~N���.�����,eX��ݤ˱�cȟ�*�׮ `þu���dk�D����B�}]k���������#V�[H�F%��߱��df�|U�6�O��4�/��Q�^8�pic0�{� =h���~�o��H�;�R
&���k�ol�֥��wb�dp7#�]݀�ݥ�y�.\}�u��h��b�u�l�.�Tؿ���c�VM����VRB��a]���/}i�d����zq���ӗS�hu��vcƔj}9sb�lK��h��r�fHw0 #׶�И�)���������9j_մ����7 �z�C�-���`<�� �G_u��&z*G��%���r,s��t&=��6���re�4^�!5(7YE���U�Jf�WҢ����l��I�|fu�`�������$���){\W_���m&�[��.�!:�4(Ͳk�a���4������&Y�\��hݨpN�[<��T6`[pe���a�e��������y4�iN8�����8xץ�o[b v��.���u%/���y�#�;\E�D%�q��UL�8�jZcL������*��@����;Mc2o� ��I׆ �H^�����@1��p;d-���G�`l<�y�xCً3=� �2�[� L�'��<�:U����(��a+��`}���d�r���a�ۿ]&V�~���^�������%��[F����p������d{���IvR�&�.j�6�դ����:���XlxVHYEB    fa00     5c0�DA8�Χ�j��������uI�^d)���b୯����*������t���(�z_*�[��ǯ&"����"X�5ڨ�^uS��<����p��k	�f�����n���G��C7NGP�8ǐ�iƧ?�ZKX�>x;˞	�d-�~�k�¤&Q�E�4��iZ5�8m���(,Ơ���ct�b{��v1;����jX�YnW��9uz�J��4�ۂ�2�U'�}K������sV��#�i�^�Ns�L������+l���H7
�j-�Q_�L|���A���G>��a�_"�̍zA�+RN�����Q]way�]k�m�����]��g]"Y��Cg>B��p�ZƔ$��<���φ�n
<�k��_�{��V�^��v������	"���M�¬�,9����a�A^��:������䎝��pB��0��'/3��QH���:��?�h�Om�@�bF$w�����{X�8�t��t�S�#����<p����J�d΅���
�Wb��Y����]�Aº��ㅠ`1��Yx��Wt�yT���9X�\�w��н�[A�o~��"���\G�T�Q��������.�3��
��bؘ�����f���8����YO�<�`Z�ŌѰ�6z��`�o��R�z�ͪ﫸�v^��OC����'<	�7�t�S�[.N�HP.�n�!���\�Z��9�X�\B��gX*E�SvP:�Y��A��2Bg%(�OĴ�#qd�6@MJa�2]5�(���'SL�R-Ju�-׿SݾO,��Ҕ�*�/�ݐ�#�,��S~e����A��<�Ȗsnv*D@����T�&�ߠƎ+}u�����芶�q��'��.�F2r
W��v�1D�ES8�͹u�Jj�A�0�j�%Q��Zj��s�zRd�T48�[�� m��f��6o����6Gܐ14�"�NGZU�9�TZq��M���FPk؉\x1)�$9�{4��у�h����a	uo P�ǵ���>���]$�6�ʏ�Y��>1���?��e���Ԕ�e� F�����D��o�1���*#aG�޺���H�G�@�w��CW��j|�sC�X0�.v���>��D��N9S_�,@�*�Ϙ�5W\�zZ�3M���"����)�x�b%��V�4Eִ�b��!���r��uSk�լ��3+��W�'J�drj�l���e�/GXƉ�/��]C~bV^�N�MRޖa�H��H��j�J/�����,:�݅��M7j�|)~�{�9.'�����,���!6u�x]����9�MUTڍH~+�a>��^�]�"��ʗ�²>�8�~�m�)���u�嵌h�h�U���S�OZ��������W�zP����}�?�9�����}<�Z�t��ϵ1)�v���>\V��ӳ�ma�0W�D�0�L�=����,8�����E�� i�F�,ī��ۏ�N�dL���\=cu(�e'XlxVHYEB    d35c     aa0�j�����?�ͬ8�^ �N���J=~Z_�����cU4|�M3�-�ӹ�vJ�L�L�z��..�$s�,8�)����r���>/��}�м�۸�ʛ6��;NA���ͭ�ӄ#i�����
O���s����0L!��m�8��`ŉPgߴ���?3`?�6g!C�-���U}'���+{�<��@S�����dKW�m�:� �7�|�H^��>MJ��Ѯ������1׏:��{`��6����ri<TS�	mBU��V�D�1l��A�~l���=��}�]�:��q�f7SڊR������^�=h��6�#�t
-^����󢶵5�$���ǀ)1��G.��-��]�R�R�'����b&�(��i�dOer2�7aT�E9�_�z)�w����7���B4~Pu$�̧��(��B��b�2n�m��iN씚hSu��t�i�G�v��ej�e�E���Wm�mD�N�*�㾽�M�-R�ܭ_����N������G��� ��௔���8�,`6T�i��Q5L����Sh��@z~Qᯂ�`\�����������,�E�\�1���C�*s�4��L�;�9���:��)[DìN�W��ܤ���jaV�l�	�����,-`���J�=� ��G*f���%������dZEr{?rt}>�`�Aݸ���D���}��	�Aǁ�.�@�A��LI o8�~,^�Q/3Z/U~���|qv�b��,iXxHt�WJh�pd�L6���E� �u��e�"�~7�k��j�l޽�3�hjƠ�%d��.�~�=+2���k��E��[�Φ�ΰ�r2��፸Q\�'�#*f���P��[��m���<8�`���'a#xr�d�תϦ���F���Һ��1)ӊ(ޫ�
o����h#XXg84�uve�d'�º?����wIw*��>/��uR��*V��4��f4�J��H�<ÆS	5�Ou���6�-SA�d?: ���g>�Bd*��]���2���/��v�U���*Tѕ�>w5�e�"��L��@�C/�/���ܞǛ��T)���М�N�n����|FχΝL��;I�v��Ѧ�i8�7�uVBw���.����1g�2$�'�4��Yf0�#[���`������r��ʢT�N2IY��X�4.��;k��Wߺ����.L`�TP-c��C6����Y��*�HM�a��n�c"�H��iI������1���g�j��K�e�)Ӹ�q���$�}4MM����?'�Qk���O��6>"C�M���׹�/�Φ��r���R�"U�����Aq��Vs5��&��Gq�ZC���8J��y30\�;<Z�SE)#C���|:�d8}��A7
*�|e�˦�W;�@�ų/�k�E���6t���T:+H�%�|�5\�?��oV�>Q��K�C�A}5�<i×��-��|a�����A߮�n(9���b��Wo�Q}�w#��w��9���W�%Om�[��ȶ���i̳� `���&�/���r6���M0�OJX���v����5�j�����b$�-T΀ON	�p5�S`�m�����~�F"�7Ң�A����\��$)[��h��	��G��%ˮ�ޘ�6_c־�Sb�� {/N���B"%*_� �h���ո�tP��]��`:b&&n�m�ppW�sǞ2t1=�*�q)C����e�^����k��UI�V��z:v�x�;A����P2�_�˄fLƳ��� ��\-���~1D#�<_�N��yxJ�{p9j���5MN=�x�p�$!�����?���@y��~F#M�+�z�h�8l�����y��?�ď�p��Ĥ���/�7g�Fv,t���]CG���L(����ը'5���j@�u��Z���̃�b��|Z�A������6�s�g/%��	:�H�X�;�N,�k��Vt4���t��	נ�siT9a���zZ�P�Q#�~,�C�a� C�6�D#�mOO�m������]P�}���LQ�"L�mG�s�E�V�k��}+6R���q$��C%�x�V~䌧np�C����(��Ȥr-�^���i�kCs���D�2�xF5��e���/,�٦����΍G�2�e�[�.Y���0�W��E{�����ger�"F�B)���0�G3��/N�\ȁ��K0;@�{�EcM��q�f��@�5w�p=:�C�2����O'FSp��ci��Z9�V0�-�-X�e��:Q�:���X^�y���Z�1i�g�D��/�)��n�����{2�N�\%�� ��&n��4a*jL�<]�GM�k:/Jg(�qC
��a�F���: D?C!�{���Z�܁��ϡ��?�9u!�E�V��j��F���UlQ��y�O�5�𻉑U���C4h�Q�P^CҚ6&�n5������7�Aѯ��Q8涝�Hʙ-I읆[��l���1	��6�&�� +���D�k��4�'��ݬ�.�JՖKY�.j��nm�!�79`�9ױ0�M�v����;����W��� �?���#����Ï����������ۗ-"��ۀ�J���"�eJ�9~M��§��!�����LϬ���챨�A�����Q�i�'A?*��&����
$���1dZ��i~ō%�i �y:fSs:��0oCk�Ǿ�����_��CaK'�<