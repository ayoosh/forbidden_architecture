XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Y`όG)��Lo1^� ��9�g=�t��pm��=��xYlw��bV"�5O��A#X�;�`oaW�n�"5��G����Ae�;�� �����P��rm����Lo����-�D%����ߤ%���N3;_;]�i�nvR�\��#�7�5��w*"��5k.�`����L�'�+@I�8{o;x}�T��d9��ϗ�t�!�N�+l�B+�r
�^)Et �	͚��%ON���zd\kqk9�Q�Yo���gH�PoS����a��7ȉڇ������F9�}�Y�"��ͳ�D5��.��ӻ�aF97*P�����E��z�M�ĉ&-���G7�qM����)�F&�֙/S�٭c/�g#�<��-0�4��tI����h�i������q9��g�����b+�AL9x�N�~\�!s�l�w#�<C�g�.�A�!��ƾ�(��rs�8'�2��8�z�ԃo�	���'�:o���)!%���/I,���O����˻ݟ��ɣp������&�ȫlIP�<�l��n8|�A��T��l��-80�&�\k�摗iBz۞TB��}�!��4��8 )���w���J<
P�]ѣ��<�ZF��s��胱��'�5�8�:wvKˣ�ݐ�d�,�>1KԌ�X���>3�`���+;$=.�z��(���2xS�Y�����n.Q��bj�,��i2^�V��{�~lÍJ����l+�V'8����L�D޽�0�4����c��(�hTw�`���Gi}K�%�R��YuJ��omXlxVHYEB    29ef     b00%V�e���qo�T�)�]KG��� z�8$��*0����.����+g�G�Ft��p�ݹ�п��"���:�je��o��'��yTU�R�j��4[�-��*_�-�X�}(��&5���yI���x@�Xa�\^�Uz���2Lب�x$�J"�u�_�����KK(�b�����^��U�A��Oת��}+��I}�g�d���x`��&�S�y��f)�C���L���N�˕T����mh��s�>���77v�k��L��:�／s{�5�/�E^����p�v灈�z����v,k++��!?�9�=�1�-rl�1�52�Ӣ`��CӘUߑ���E��4�m���j����I<�6�a��B�R2�D�Y��p@�"Ů�.�6�\--��E�(�]X���PY3ҳQ�} �j����V�%#��B�g|�⽵�}���TL�s�{�$�f���$�J����F�$:�//ʃP��P&��Ub��������No�@��h���|9ig�B�^G0I�SNL� ���yWAQ��_��^�21�Y�d�s�b�-?��_&�<t�/7���X����nҲeJ�"�0��P�ib]��-|d�Ȩtu<��]����2�&������3�pW�(Rv��e�?[�4$)Ơ��	�>d��N[�M7���E�1|��\N�ZϢmo���f�JX뫝H�eF���J����U�`|B(��I�3 Hf�lI+G�4H�z�q�a�A����mG4���z�ۂSLH�6e��O����i��7;���H�*�������Yh���A�OV��ɑ_�%q�Y%@b+��AƠa���
M�Q�l���Y4�RM�fW�[���J�U�k]NzW�K�:9���x��rw*rTK��XM�V��+_����q�h�(��'��M��1p�O�ؘ��/�b�� ���q����!��,.&
��?+����d�7�`7�I�WE�s� ���L)dO9Z5N�<DU������A�il�Y˺ \
s�r��N����{Lg��cs�������6�׶N$�Ĭ�A�)z`ɞ�'\fz$''*ܝ�=z:�9���H��[�y��?�sB�._��u��Рoq�j1aZ'b{�L	g ���1A�8O��W%��JVYJ�o�Td]��q���H?�̞}�G�v���e�F!�ԁ�.�-����p� @�N��V �L��XP-�41��Ɓ�*�j7ؿps�*�|��i�|]��;��#����V���ρff����W��P�*������y<Sp�
��]��P� 5��ҀO�˝A��9�sܜd����(]->*mP���v�%�X��fS"�j
�]V	B��LJ�"�J�<����h�R ��-e0�Jpͩ�W+��v��K����(Qk�f΍,��o{�@ ��/nq�31�,-M+%�t
�3O�IM���´�������t܄E����fb�!�0y޺nëo�nmvG&�eu�U�*A�M��x	�����	W�&ϰj������� Xj���Z�8	���wO(�O�P�x�D�>J,�'P�̶V�Cd��Gy�.�����8�g��9�J�`?�:�6���=WtI�l�K�౎���ud�a�4,Þy��i�g>�Q6:� �I}��0�>���HC�"'����(6xG�$xx|(�Q�X�!��I��f���W��w�����i<��E��!R<W1���뙔ڝ�T�ʋo8�?Tð+�P��'��z�i���&�8DT)e�r����;�����w�s�P�.��7�T��ϸ�Q�0�T�;=����K�����}��*�;=���ϼ�C�4V1%�/y����k���,P�׮LO�^&�$=yٱn5�G���ʔ�=����]舋�\V�����8�at�@�����vZd))��5t���+	�=����(����:�;b9�7xke����B�X������z������}�P�k�ۣ��T����c�sMy ��]Ď��m�Q�&�-�C3[���މM��}� Qm��aL#�%E�XIy_h�!>$1�m!�
V~*���R֌5*�*�X(��o��NexΎ�Vo���U�`j�R�fR�TU�%˜2 g�Gǐ����p�(鞍��}����#����z���9��ҷ�(ZEBʣaI1O��z �v�?�+ڍ���}��eءԹw٥D[V̽T�>}��笾�mS~.�fyK����(Ԓ-/�9hrS$��vn�|ا9�a� 8���J��4�1M3Pe�(X��ݑ���&U:;�7^m�4�/p���DbK�k���Y��P��UMɞ��*��^�k8�`;�_�C�#0��BD�O��.)��D�_������b�sbߡ�����8sz���wB�Xi8�GEȕ34�;����0rZ�
<�`��^���I����5\ID�s�	��>&4����r;�mC��ݞ��w.$�*ۇ$�?��r��fxkt�&j�?.�h? c@r�h���&�AV1�wΐ���)��p�	�Z"��7I�%��鷺����OՓ-U@�lU:y�4�s�)��܊X�@_�ļO�R��2�R�'1ψ̬j��=�$Xo� �&�T�T����z/ ��'Ҷc�m��/�N/���uݵ^S[�/0V�R�6�7�V���v_�&�jC�zn�z��^�.K:���Z���_��^��먳�i<\	�X��5i��u� �M�מCK���i�; I\q���Q�� R�t�K�D!��������U�[ԨZ�ƈk