XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����*�_Qz�1l�u��V���9��]6b�֏;���R�#���۬M��[
�Wp�͛N�	������+���M��7<����E�����=!�� �ȼ�uϵ��g("�.z�.��A�ǘ�x�ƪ��|/\�u�v`g�D�dR����#f��m��m9nt�%y:u@s�+�m@��g����f�l���g|T���X�h����F��X�p�ٝ�c�&�}�8V�}�2�Z�k�$�ivJ"=��8����*xTh�܊��{S����m��A�ʻ���U�`p!���1��?u��� ��^]�6o@��K�O��44&���y����3U�)��I_"�plU�:z0�kb�j/��]��XW;����f�DZnkL�c��)�٤hA}���.P�|�f�+6�S����|.�!{���x�O5m|����g�N�� Y��I��o��)E�-ҿ��D ��r\4�5
.\�}ާ�\�|�w�]������DǇ2�Lq�ɕ�D2ˠ.�
�b'hb���
�D1��(��q�݇@��{4	���9�J���/p���]�"�+�������!�O"w�����N��g��Ђ�(�?��ƟAL���<Km��%^����5��%��/s
��C��b�X��g�eq�6i�j¨��>Cʣ�����))�#�@ v}��@��G	?ɔ� ���I��	�З��0�����$���	��@�|#�_��;��0Nv?������Y~�߮ӓY�XlxVHYEB    c763    2600�Z�"�W�^�զa���b��]��~k�=! �ݸ���^k�1�p�b���O ẙ�(WC3�UE���|�P�4�cW ��{$�߇2����L��{��!$��R� ��:U|;H����Ϥ�ږ�Q_����h�
���5�3R���EP�����7~��jvڡUe�M&�ظv�y��d-52�mn{G�O?���Y��S7�/��Q���S')^]�ޱ��y�̢���I�[_���@��~Y��oW720pǤ�I�V9*��%i*��i����ƈ'���[~�Y�`�j<��hy/S����e��?j������AK�i���z�n=�)6��SwщxN��N���T��8kq�����*�8}���z:Q��膚y�@_�_t>;!��:_l���v��ɥ �7'�l�4� DY��ҫ�q㹺J��y��(��pD�H]9#��u5X��{D��=C�q#]�B���1Q�>�fRJ>Yv1 ���*�?�{9`N��.�R�S]���v�����FXT�th�������T���ݰ��Q��\����Gǁ�����f0����2F��I���M�"h��l�nuD��ϒ�2_h�r]'�XU"�Y$���Ƨ�= �j�a���ub��+ܺ�w�o�ԹO4�;�(��S��ޘt]`jN��[��W�����b�[.�aA�(����0��^��w�N��L���
���[0����mʌ�jc	�wv`2I<��H���4�����j��RA�*�_D�_3��M;5���@m�I���Ŗ���k��G.V���=�d��6�x���+ѥ6=&#��J1n��<�%e!�nɺ���ħ'v�*V�>t/�#��-jḳ ���6�ߌ�7�Ϝ={$X�AltI�o���_\�U�c�#@+v�h��YG�P�Q�h�F���#E;��^^����#�O-�Rʎ�3�wAY�b��$��E�nB�0.m�#s����D���&GX����྽K����`Ө��)8����:�w�Z1DV%���D�����`�*�)�>����4T���������3h�a��M-߿��\k�[n�_�ҕ�6�e|��H���Ǭ=u!�3f%�}fg�`��x�L�(K�c�bOa5�.��%��ވ�F� H��!bԯ�H�at���4>s���a_`�Յo���T��&�9M;�J	�)B$aROQs<�Ĕ�/��㚜�-2�j�r{G�r��� ��!	)�_U��Ӎy<��p�eP�qlr��o�fP�<�w2��wp���4S���� �%A>CH8xc��1����v�l��:��Q\�]aM'��Am�l��]��|����C���f�ߪ�!H(���C����qr���u����;ʋ���Ss��`��nĎ�b�*]h#���
	^c��Q��o�,j�&1�nӮ.����Ia�*^6��;#G�8B�O2�\�uh�m��ihBl�o�����;��,�@�)��/��\��f��t�/E��u�]�#ǀLI� �1������q8u��'�@��lZ�*���Q�#̑5 �����ωQq��V7�4����fy���j�c�I���^�|��J�i+Hg�]�tb���~D�D^�����,�z�h���V�$^�iY�����]�T��(D���wWf� �^�O%)wI����[Qug��.�,OŁ3�K���� ��^�kf[�]{: g0�c�K�Y�E����I;%ֵ
KU)����/�h��9�7��	_R)��r1QYɆj�;��Bk{�H��]�
���v�A���e ���o�!�1����0�~�t�z��UJ)]�q�Ͱ�m<�C��C�2�)c\3&e$x�/Zh���0jV`��qV����[Hb���\淘"sJ���*	�%9CG�"w\��,-��� �H�����ژ�2u���s�3@����0�EM���κ ��Pŭ�u��k;�{�(���ӍE�;�kw��|}E�?`'���,ǔ6)ˣ�{��J�{+U'v(!��4W�r\eu��Hm l���P���q٩�|#\j�ԓ�0e����qf�  눑�|�������yviGXU�j�x�ЦL�4�lĀuۅإ���ί�m�)E���_g���ky�I��ML��̫步�T���� �f'���(:�`�
��C٨�˙M��̏�ۖƮ��r:Y�?�W��Z�E���nayދ�RSS(eP^M��m�l��C�j���mG�b�,�.�@�K����VDj�p����lD�أsC���x�U���>��T�\r7�U������=f��u&1Ϗ���i)�4c�D��ʠ0�
����'�Q��w"w���l�皦hbX�X&ǩ'�rlh�YbV�񳱴�A���{}�Q���)A���<�Qg�	�p�Z�v�a�mZ_y`�s@#���j�.a��}��;9�.��R_��>�j
���d4�O)X�W^�0=~g-/��L�4���<��-�lWyz	� GEO%$ǳ2&2.[�85�vZSfQn��f�:�YB�&>o���- ��|�}X���w��;�� �fqX>��Oޒ�i�C�/Q�+ZX��a�g���;����F/_R�L�� �o���
E�J���&t<�9��k�F�x�-$s�L��8?돛��$��(���j-�M9Wg�*>Ҙ��n6�vE=f�A!T���������1�  U�v6����z��K���}�a�5>����'q�N��P�� -�#�aw�}���[���l˙B��d@V����Zޝ����~����O�{���'��%�1��@C5w�����=z��fC�.�hW*�0ȜɃ��}�2��y�or��eJ�Vr}:OzT�=D�t}\!�B�h�_�ԨW+b�@Kϕ�s贚��{��	Μg���s"���#KO?���9H}��c�&�f�U$�BP���c_it��j�ӱ�r�<�"��P�R%��L����M�ކ)��}�LR:���߅��sqo����<�C��f��r�}��z[�[p����!�3S�6J���~(�06�ɔ�ս �7�D\u���J��)�t��<9���V?���ݲ�ZW�ڃ���@:���ꁐk������c�.J���)��:b\�S�4{�P�v���~+A��r��k
��|�/X��d��$D�o<�vM��Q= F�</k(�A��2��1�aX7��z��3�rzp�F2��]Z�<�q�QO⁆E��#��ƄJ�E	:V�e�����BZ��H�ds*�m�/M�����! 7�V~�h��͔��+�8��(��%N�D��Ū|'L�nI���N䴉oD�_&=��jg�"��kO<�H�N'�-�ׯ�Vbsp�����C��kmx��<�_c�ϱ$s�bު��\\���#i�M�Gn*�x?������rZ����yDcM6@`s���q2e�� KhK��(�<9��Q�hc-kе�ClP�����K�Z/�����b�g3�����+�U�$C%��U��I�)�"-���Ŀe˓��/�aѨZ��o0��C�%˸�7���O�W]��q�����y���ǂf�5���l�C�*SS�(lC���uǫ����������,�0ՏAc-G��	����M��s�3 맆S���.y�I�����K�?$���~=x*N��dwOi@�wYbf!D��!6xE�Vq�%C�	�� �l�b�(�������[z���a"O%ͤT�Eb�h>.A�"�9�%���}�$�S¸����wJ<�Z�����✞`��b*��n���l	���^��#��ϱ�Qt��~g�3_\����j;�xyd�݁� ���!����]���+�P��t�4�����32�
[uI�f���ąP �R��_8�*��#�F>��u[�xYe*@n�4� ���⃎vT)���R�p"������|{6���3F-�{�'`n�Y��݁���h�Y'U�P���K������c"W��7�.��L��w)I?�)�C-U�1��p$����77&S�U��Ƅ<����@����Ո�t_�&�}�sB��O��~�,�2�BL�J�?�'t!�Cϲ7�WK�~Ma�T���$�]&&&F��b��ش�|�Gg�a�=#,L����0∾��v�=Bk���=h؇�x3X{/��#U�o�T&)̫�/�4B�}]@��\P��)Y�*���ui��3!��}�9�K÷2ς)GW�D��\�f���x����lb�͌��_�Q]L�����ڧ�֫�5#�[h �&���"M@�SumC�y������0�%���n�TV����;j�ϳs�P��ѡ*6�#��0���vj�m]�Xw�߫�����8�R�����6? �Űs���)F��O���§*�lI�j�G�*�#'|9�����k�'����J��d�0οע�l]zتv���h-睇�~d�&�0��H��Ls�,��� ���M��t��k��Bf�GK?���+|��j�lH�r�$D[�{B��u�˕�-�b���[���z�D�˔�����E��\ĺ�o|j��,@���Y�g!��}Z0"��q�y�fT�@u�p�Ig�}�ܬy2V���#3�G:��H$��l� ��u�aL�~	�WQ�&���3%�3ތ��6��[u�E��זP1������8�
�)��+�������I���+��g�z ���	 ('�zߓ~���]i��V����-�&Mh-@�g}2�v�bҳ	 �:��Ux��B��(�Eh<���אVS�}�R��J�KM��v�X�]���kHg��E*�X	TE�'[!xĒ�T�)��
���]b���Ċi�0��K�4��|'j>
��n�Olg>����_��V�%�.M�34 �^��]�#xv���=)n��,����'�O�ee�l�:�v�u����c��>;v
ݔ�T�9&0^:q�������;�e��-�b��E�B��˘�5D��1�8�ߖ�%����y�Ś�;lN����|����/�����}Y�b_	����|8_3�Y���<�s��mzR߱<�7M���g;�IT��%�/R/W&�Dy�L�F�+��݈_���F�(�u�%���8������H��=��]qg;t%�'�X���/me�%>�ݻ o��>�|xm�)��*��8	
 ���p�<�s?eC�(��j���o>L�{ũC��* ��eq�f�$�g6�V�_{[9>��f��X�� 
�'���8�f�z�:�=`�OQ�X�o��d?��SÉ��2A�2g��{a�W� �������$f��eSlZZ���j��=G5�5����h�;A�5J�o�PY�i�ޗ��4^$f�%�pq��D��{��e�mvx���V�c<���Idߑ�Q
��|+��)�u_��,`�%Ar��< po�{�j�Ѿ�3Q.;,��M��-I'��Ɂ�
mA|��1i�K�
�	Mj��тkoI%mo�뜰�޾ S��������w�2*X\%��������Xň���l���Q{#���r���K�{"��-��L�U8p/[����>⪅�}���#Ǹ���n�I���^6�Ų��33ŴOD#��2��6�&�L���j��G��²��5�a�ot��7�����e��H5�g.Q@��?�^�,��
'�(���/�#����43û�~L������+m6q����{F#^�ۼH���֎�/$���K�p5<�~!�ɩ4�_�j#�u�X�J�j:g�:5�;0�9�L�Ncf�6�>/��������	s����w-��'T�,�^	����B�	{��>4N�^���g�3��(�E�$�8}��Z>7���;$��/��oN+ REGMY<����Ugi�I����U/7�Ʋ����8��SE�$�=V˖���b���J�Sgr_��������}x�n��Mn��0/���DY(��hO��J�!�4e��"�rp�O��v���,�'��2*^=�@mx \���b�=��M�t�5�3�}�tRO�ό)w�t&T�����&�L�V�xmK�Ϗ�̄�Z�kDJ�N'	Ư�4��s�TX�4gP�1A�g�j�4}��t�Cf	8�����C$CV�
=ߚ����w�[��=�แv�< bv���e1�8r�姷�%�7sS%F�iԋ��u7��*~�J���7�ޟ-fC�����"OR������u)�u�CJ��M��$6��o�srjQ�Ԅ��EQd��+;K9D�K�K 퍦���������l�bI���&<�(h�5��1�(��τ�_5��Z_?A"�E�+�]k��c�P��������x�F�5vT�����>S����q�jCv���渡2Gi����. �������E��?�EŒ2[��A���� CZ�Jð�i\	��0Ya�.��;�@|��N��+y��j�j���h�9�<3پ|�b�Qb��S���*9�rM}��B�曒�MN�QՂ���E�h*^N88	=�2�M.����	�E��%�~��Ӳ�ײQNp(G&G��V9�A�ӱ�8��A��f/�h���(���Uz��T���Q6)�f��{�YC��6�2(�zlA�`�m�j2'ǚ�5UuAg�$M�	��sƐ|b}�Rj�.a>��.GC��Q?�i���筪6����'eC3Q[��h@�Z���]e�R�Wn��qX25}�3_&j �7��et�^�S�n踗[G3B�~�[��߬z�X� �9��H�`���%����+-�sΦc�I�:�� ]ͽ��m6��2��	�xr�,���A���P ��k&r�@�%|O�[� MF��]�Ԥѕo¶ofZWH�p65�s�9��|�p��� �e��܇�E�t��4��;���m�O�@J�c�Kۮ��s�kd��b�y�q����Na�b�S�:�W�^�l��q,aa��s�5_�[�L���w��R$6��Y�����!;x��N�|G&���0�ԼW������K����|���|6�"����y�;R7.~г���<|<T��H��d�a�@;Az����n.����8~s���uQ���ܟ7�[���e��������A��Y��(ı)8�����k�W?c'�ғ���(eWQ��cn%R	�ױ�H��T-(4-�a熶UN�ӈ�ᰫ�V�,
7�n��Y�׮n*��	o�(�#ϨPR����ي����^���@�\7�ր�9�f�C�o�L�HeZ����VOd�B�yĝr�$��>��$`֔������8����$e�WBa��t� ✾c+U���R*�bA���Q�kg)������RךC�6זdH@οjl~���[��߀��7*!��/���w��-�L3y�����/���#fV2�eqr�K��p韅����[��KV�o����x�t{�¼^RyT�U��Ko���V�F�L�ƴ�ծ~����mB�|]�Nf�&�0+}��K���Dk�-$)fj��� 2&u|�h�|�xa,K�g��<^�S�� ����k`�c�#���81�o�V�G� ��=��S.Ŝk�YN�S���TN��2Iؤ���8�!�����ɔ�}�\!�Z��,���w�(OT���la~\�v�q��2`�����=�%�IU��C��Ƃ�"6�4�������6��|~�ѝ(r��/�������� ����7�b����[�����n�!��ж�^�G��T*ƣڅ��|�P��u�c$K�]�g�����~cݪ9:PF\�=Vrߠ.��rġj��Y0FI��8��ܾ޺b�Y�����օ�S�]��|w\�<�x+��C�_���I|t��Qcp:;ivV�,~�6 �o�����\^{��cɜ����E.�J�(�ϴ��S�-|.��YeC��5��넙��Ŝ��a��"{	�c�6t��瞦8�'ëQM����>�;�lyJf[��s������#�%;m_Gg�㲝J)pu��`8k���n�I�A'5{�s�x�vY���»�=���~����~���wE�8�؅b�y����b��q|hu}�&D�]U�'e :�g�v����7�s�U�*�^��
�8�C�Wi�DT��B�:<.eF�=�Ƒ��2P� B�@��YР�/&?ۗ��G���d�E)ӡ鵒@� ��^�+gLi4����L��vV�書�Ӛ��n�o4ڨq*�X��s�o<�j�d��8�?p"p6%���0	~��M�3��;xEd���B�H۸"�=����)�%xbB�B�aO��a��p�a-�h�sQ��ݢ
�9D_�5�c�����C>z����cnqk�A�� �Kk�;ui��sg"\�씣o��Z��fҕ�x']$�]:��Gs�є��Xjs�c�J@�q�;���/�CK������ō�P1H��� ����ʘ�_�������73 p�(�`:�v?nxn�#1%"zg}jmŊM���гa�\���>���+j�%[	~�_I6���Ѳ�վ�u���>��u��3�D�;������u"�!+DR��[k闝�ˊO�m�E��^ �0Ӱ`g�?(v��K��r���#B��m��Q�I7*׳\%��2��3��X	�s�SUv��PU��Rk�@�ڡ���ӕ{}��" 7�3�ן2Okg��X
���o���[����B�&L�]�+���N��t;���y��k+�n<�ͮz�3o)�W�i����a�})$9�C� 9>
����R�k�9��Yӹs��~7���x������{&����E8¶(d��n��||�Ƣ��*��S���=�Xw#�V����M����.���n�l��&*�t>�yD#��>Ȥ�;�޲�j|}>?��P���mry�����Q_�ةH�aԦS��M�)�ek-�|�c�Q��s�z<�x�Шj3�.����$\��ף�e� �Y��#���{�l��J�J����,��5��O������ >��L�i�*B%B� J�	�~W��0 �sf� D��Y�6?����H�&󿄋�J��g�[2F��c�6I/�<����z{C��^���i `2]A�plex]Y�ܚ�x.��h+|�r�k:=5�`.O�����ܭn'eG�4*(Ha�"��)�í^v��L$�o�h�d�~�n�-���%���v\���q����ʈf�X�B�x�L��hD!9�:��q�Sy��{�xy�6�̈́ƚ�A�M�_O|#�RZ�M�l�dVm��̺�#Ѷ�H�]i��wt�R-���m�����ѩ��^��9�N.GL�_j�ݟ�F�Q�]ԉ����U�Fã[���l,�x4�a= �/Vϫ����L���L���]Jd��\>�bkl�������Gr����I�pu�d�����]}]z�*H���I@�VWsY�L����r��@�΢�����m�5�	'��^��sd#ۉ��C���,`���T��� >]�f,��++3η���=.Wٖku"�M%I��)xI��~��좾��	�@��U���ZC�P?We�U6b��z�u