XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9L̓t���8�W) m�"��V�O�/C�8���3�pf��']��ad,�(�GwiK0���Q��~i���К�j����P|)�1�:g���U���к�Q����e)���|��N�G�F�:M,6W��\�Y�o�.�W��j���xZ�ԗ�&���[���쉷_�h;��ˈ��{Y����#��׋�|��(���Sk�HNQx�3z���lLo�?s� Ϣ����t���p�WrWcH�|�ZkѾ�>�@�v��r�DJ�P�+u��c,��z0Z�$s���sZ��?�	��33�I���+޵@.6a�Y�K=N����J�����$y�\�.��;�1|gf�}d�ԧ�P�G�B����jh�7�H��n�e��\F}��<9E�a���uR��e�K��U]���
�Z,v�/��T#�ndH�h|s�@�V�O�ɏ_nS�Nh-*$��al�~OnvlH_����|@<���Cq��'ߥy��\0$e�O!�q,�%s;�)��p4�l��\�u�3<�߁:vĚ��>͗�,W;���1�᧟0�P	EX�!�5:q�茄���56B���0�?����D%�`��|C�`E+��g�0ωm9h�C��}�z����b���Y�,3E� ��ެ���$J�D �x��ͩ������._��1o���m�y����$�-���f���	I�N��f�ے	>�G��|����)"��H�JǺ�yf
��,oD�O�FO�:��z�� �jW҇XlxVHYEB    fa00    2470{�Z�%T���}����6��Q���d��]%W�;7����Tu���t8h@-q݌�9�O�G�����h'���|���,�RQs1ZD� U�L�����`au�As�<�+6aT����`�~3�ę�O�"N��(�oeS�'�p�X��<fr�S������E�d��a39IB�`����L��YTjZ�c���
��~�ΩD��A���[5鍍_,w�������ȝJj����7���r/����l���>��$���$�-�dR|
S��X�f�$��0�F�zEn�f#5��_.�6��/�'l�K*|@�F_;;qe�g�i)5H�x���y�����6A ��^ q"���r)t(��{Lq����X��^
W�.��һ���L��� |^#{�o`�r\D���Olg�d��|��D�����!7Y� ���P9#(B�u{��"��l����JB�ݢ]�N�� �4����A	@��D$`����{���_`���!��D�w�XJcՀ;y�	�WS�K��ȍ��
��	AH�R�^��*�9���^OV�s2��78퉟)�:��O�Gbs�^��P�&�Ww�� eǕUY�$aְ�!���9�Z9a�Ə�����xO����oIY "���dyÆ��M�LDky�xF�ֶ�������Hr����Z�i�M#���4��nv,)��ϥ*w�1��=���ѿ:k�ޡ%��X��<��7΂��zO���n�w�hʪ@��nH��o�uP?T�����63��)�D�����)��*�ܦ�e��B�'�3	ۀI��7V���-�q��=�����_���&�^غ:@�x���$�ω1S��BE��L+��,f⡐�o�	���9���ऩ�~�2���JR�]7T�;�+<m|G��Ѱ�\��igOVV~^�Gqï��=�ҤA���ܾ2���Jf��Ce�T��|$��g����ӄ�����~�(����L��μ	�T��Ei�|��c���`L��1��11�z1ƇOTv�f��Na.�l�}��5�����<<�RD�~�#�>��&R���j�e��PM�E4�u�$"\��oZܔe�&�v�UX"���f+}ֿ�����΂7�2�=����Ο�V#�s
<�ռ��Ebo=/�ͽ!e��R;����[+n}%��]���$�x)=k��[ߍ2e���C��wiM��%{p��� �I���q�,��.Q��맆D����7��嵆���Bim�H�֟UTñ��є��`n]�A�!����ZĦ2E�ݤڸ@���3��.�5j�!|{ή�<�Wp}/�R�1Һ��";����(�B�@sUĩ��o!8^q�	<swZ�g����y]��JO����C���kG=V���*is�~z�_�M�'[�>g� h�)E~���Y���J~������BCI���w}��4$���4�[�?�m�1Ъ��#��uK~d���r�����B9��$\R���c,��nQ*v}���j~FH�v�G�����7�`QA��dc��p��^[A��K��X��;�C)Y���*Ɲ.��ߤs:]����e�jw�o_G�~��E���SI�N!Q��^�1����;N�r\Mk	GPo��3��,�(�ڶ�0�u��h�HG���b%;'��9,)u.�C|�`��_�]@L�	��A��3�)�3�G�Y?�[!��[rm�|b����'M�y
��҈.+�rZ�н��o/�L ��r�|6����y��O�������Y���X��*��\�="�����Wew$� �/��ض�/R+4{ɭ>�յ옠�ړ�ML���2��sI��?�����)c1ӼY�v2�`̨S��!��Z]��X#܆bY������#I6�ޟԧ���\��|K���U^ ЍS�> :��mg$�Y.�~����M��hЧ2���#��C[h���YK��r�+�!b�i����(�%C�X�X#����*�ԧ-��[�o	g{[�}���e�KG/��Hs��a�r�Ғ��7���/2l���df�U�/���H���M���]��Е��X��Ah]��_Y[�4`?�f���ZZǢ����7F�:5�M]�A�=���c!(�6Y�kK��P���Nhմ������
:ޗ5(�pe>�
I���r��ǭ�S>��d��
�Q@�/ �ם�T*�3z\�<gq�[�d�Z{&$h��EM��v�(3�̌(�ie~�'����~w�*ɺ̳�P��Ix�����Z����&%����W� ,8� &2T����3�D ���4�[�:�X��:X%��3��V< )�V�%��W�OT�"5SS�=L�>�����F
�F�&&at�9$y���:hh2!��ga̢O�@���iC��y�E[��	�;a�i�&Ķr��q��h(�Y�˅���Δ�&T����T�ƏHqq�Y~�Z��b\�]!�HٞIT����+�(aL�S���eoL7#�\�l1(�q���V^͗TT�원�����^`�ﲇ�6x���H{��$�ztݙ��q3�&�Hw�9c��s��T(�����~vv�n<�.���Y�-y���!g稄@!��ww������q�5���M^��|Jʇ�^�8U�x��˥~1�v����ǔ*�5_cV��b�f�b^W������Cf�|}Ǘ~�l�Ց�0z(�h��V)�z��Li�kf��_�b��ܨ�r�T�׺���=��O�:?9X�D�/��\8Y��^�UŅش	Mb���<
Ң�,Ӡ�?H&�u4�rO��z���#CW�/�F�F��GqSuGkl��� !P[�n�Q.���)י�3��+	!�l�v�>&c�C���^�i���捛�)s=(�S!	�.j���^�h�>7�Z�a�1{��)��Okߏg���$����P�\6�r�Z����ƨ��M6�W���)V��и1�):����y������WNl��w��Ɓ�{x���?D��]�	��xA,pp��g�m�X#��	���a_3�_4�+/�pO�K�ӭH�f7ǿ͵��oz<�>���g�'iY GeYXq��ݠ�~���`������P���@)��^CP�Ai�0�]���:B��E��"�� �
�@y8W���G����a��M��"B3�������)sX��)��T�"��a%�G�А�6�h]�( (J�D~J�v{��1����t.����]4�F��k �f�9K���xTsI̝��l���3�7ֱ�L.!w�GY_j��"O�cc虰^F2�'�J�����b�Su�y|�*�mw�r�y8
8���JR�(q��q{:�wղ4$��|RBÂ��G���vܙ��]�T,fH�O���s�ce;��Sp�/�y.��տd��'�G���d(y�qt` E�7�F`���-���x��cz,���da��X�]:���&�����"}����{+�������!�k_����ve3��J�F������Ѱs��X�&"ݫ�w"���0�R�? )�R�;esc_ ����
:�q*@ݢU�0�1���y镙tm��ơ���Ύ4����$r�=JL��:)��$�Gn���<�V�k�Y�c3d|�����?k�R�l�5���6��`$��-��9�/|.��uy8+�R�Į��b����k�}Ў�cߓ�4^����HzXI$�݇�~�p�4�ɕc0�14�����휦J��qm.�����k�kVs�XQ�6��%&�� uo�=����0�����b@�����Ƥu�u#�+C2ߟy�G���0*����d���O�L��J��J>6�J�P ��,��g�bR��XC5	�ABV�z�2'q�N�����7�ҦZ�@��|?6?[߳.��1/�������� �˶�Y�t�*�wwN8���^�ixN�GN�݃w�|���;��OX�{�F2~k}��Bi�C��[��ձ�{�zqzp�]���C�j#���$�b(���3K2�e!�)��e#�h������$y��#z|����^G� 1l��e�m8Yr�q���Q�6��A,� �S���g�� F\�fiD�}�N,+,�s�ȑ��%��P��ί׹�"�Fj^���k���
2�zw���)��KX׵ک��zG�W*vcY7��kʁ��f��4��sʿB6H����妡��׺�>f��ɕQhW����k�n��|�b�P���X��&w�%��?W�H	��?v�"j����}�])��j�)�ђ������sLP]�v}
��"� p��#�:�s%R��
��x��;��]�X*��Z���S��U�H7���m��5�W8w	-|F��@Ih���{S���r%�%0��t���w�S���[�|��xx�d�5臻Z6�v'����m9�����O��
~Oe}IV����cI��i��m��(K[��5/�aa�0'�~�;���9�0 ;�
4Ĉ�`h���ǎ����$H8��v���VJ�r-��aON=�Ao(��;~������l�K�o�/�}�c*79S�*m{���Ky�r�󽰌d�8���`����]!\0Hi=����b�o	�ˤ�=����4�a�0�O�2�z�{��KR^W%�F���H�ѝW�9j��_��8��i(���)�I{��{�IЃpr\�'����(�������ǔ��HQ1A#�%�Pu��O4�aYM��ݹ�޶�j�[�<F��g &�
o�Y����Иo��n~�y"����L�Jɕзz�:;���gB~
MdӃ��g�.*em�U���9{T����D97��,���0OVcJ�����B��WF(f��)u��L��흁�:���{��/
������[��h���cB�=�����!I�:L��U��x���p���K�t�����,h`(�:<\���hٟO�3�����-8����Iv�Oĉo��n	1���/IA�y��%����eeP��G����&�iӢ��]Z1I�R��W�_�_25�)��v웡#����2�`;~|��/�򿷗 Q�U61`g�8�Ɨ�eBj�ZE�k����&,����9��PP��'��9,Z��1�`M��+_e�>H>������^\���/���<��!Ɓ2����J��}6�&��P�t��2:���0���a�?6�G47�x�X�Ge���� 
��;���{�dv�Nq��i�O��P�{�	�,�̘�죍D��G�F �kh*Tl01qp?������_�V�P�64���ݠ����9��p�5@C�����:B�GI�L���j/^�����&���^��j�T[���Գ���������V�t��t�"����}Q4#/�hڑ"���d�@�"��ˉa�����&"��@ԛ�3�nV��BJ��Q~ȵ����#��R��+���>Eo�}�����ˀ�LD��w�6���o�d���O�m�;�vT�z�~��}�ɕ@
-�m��ƃsĻ�c�>u1��~Q�oD��~L�Ж
< ���<'#�S�f�0W���	�0�{�$�q|[��p��(�Kc�
r��g�t>�\e��J@�^Uǉ��`�	�LnC?�^W��E��s���v��9��]��J,5�㫐�{g����Y�::G�8Q^rg�^��-�C�my�Hۛ/�&��Ռ�V^�K�K-A�ˉo
�FJ(�����D���f8M}dA�u�Z�X��ԝCZLPԓi�Y�U�F̂����{���x�h87�\/G�M�������TYsǙ���wg)m�8g�c�/k}�e�:/`�Wе���73'0¬������{wW�d��LI6g�^�V��l҈�rK����}?��UYi��rKZ�)^U�i<.b��ԛ��@��������F��Jv5�6��ii,�L�E������oK+C��v3W����]A�E����)��U
��ܟ����t3Gr�M�8I;�/֐nڼ�c�d>�-��Ȗ�AF7�����O��+�
Dލ/�ɘ�>h�9pDSV�O�|{|t�q���]6���(7��on���h\SL!�|��G�0(�[�b>����.�й(�C�&�� ssI�@)��Ŷ}���u��o�0���qBL8�N�勮u��Դ�L7/{\�>.�BB^3�D�r���04�oe6J��)��G�ê��[��-C>݂%,A�>O��i�W�!ǰ�H�;@��$i���
��C���J�����P���7�R*
��t�Ci��`� _,6S�en_�	'��KHIC7H��Iٸ���C' <�]G�"����>Ɩ�9[���v�A�`�����.�Bזk�"f*��m�!~�����Pp�,{�آ�e��ïT��u�m�R݈,p��Y$R�m�i�Լ\l�ydUm��<�
-�Y-�a����$�W������/�A5+��Z+����k�
p]�K�=)fCO�͟�6� �WF���AS��Y�e�O�u�)�{�&r�;')����E�:[��H+y� %�b#�]Rb����p�օV�<�!�S���}���,���%���R%�Bx�?�U
��f����:D�������	�f�h�=���e��,#:���h�
9,k%�A���h]�����j$F�Y}��W�`v�t:6;<E�uM�,�MOq&�A��O	g)WOo�tewtZ�r����>q_)o�ك`�Q���&|o��œv­�G�ڵ�ī��n5�c�Y�@\���~3��uh�Wl��5���t_�����*�)WǶ�?��F�X�<,> ��q�k"��������^L�����Aٟ�|oF�	���k��b���S9��y���C+R,F��+ ����TY�|V]�v�giu����ܯ҅&�>}D�d���e�Sq|�z"�@K6�3��Xb>��;�]ܷ��tũ��E'��W�TS",�m ��E��U?�ry��9�ho���	��%/Y���؝G�tMHO^l�|︺Bv�º��4���q�	�|G.g�z;H$��c�?=�H��G#��a�=���<1�8�WF����ԕ��"K8���vb|Z'�n���î|��+o����B��xr���	U6@e�c7������~>dc]�豃�,�IV�d� JB��pS�b�j�\�v��4|����{-�����%:׶V �bSlR�Y ��y��LC�+w.f�RC?��y ��n������Y��}�?g��d`��=���(��<�h�ԛ�M#xd�h]L���>��R1�6�)�ؚ����.Md��T�K���I.�k�>ljɚ,���v(��	�e�����Bm��9FYB��W+d������s���
���o�����+�̆�?9�cKr�l�إ��K�����kH\a0�~)��kU��j["�3T!v.�zЁ���(���Q(Y�"	��R~5*�{|i!�����}�~���D�?�5m� u�<��薦�ݿyS2��<��NҊK�MW�U���%G&�v�K�|�������E�6"�&r�W��n�*��������D�ӄ��)�E�闸`��46�P_�>����v5����M���k��mR$ZƳ�����F��R@�f��@f�ۙ���wj�14�h�KZ�<[����-w2�n�}�pأ[+�[?5Ľ6�{�u둁��1w��꜉�f����mr;Uz��b���Ũ�Dhz��/j��XX������$d~j�;�^�������\)��8�!who���3b8�:X1vm��@]�W�z�I���FR��bG���Rر��,�f���H��?�l͂`�i?��e�����e�����5.ƚN�{�{_��5}a��O�ܵcq��F0ZX���6��������󓑟 �>/�M6U��d�G3�T<f�Fd�yF�ɳ�5�0��l-:lW�ᚕ���>��H1/��3�����5;��l��s�6H:�)��+R�ɳ������?O_��5i����2�#���;��n�N��`��GҀ����O�C	tÚೌ�5^��k#t|���j�=7��#�R_Hݰ���p���?�Jҝ�R�㰽u��Ȳ;�L���g�y�L�8Z����\I>wQ���/)\/��]@~s4?'&Q����(+��(�$�g{;{�^Qr��>^nߒC/�й]R��x���a�����c1������}N����:�\�#��..&�,�����Ctܕ�\��Z�K�D�G�A�K���_�����a��^���ʥݭ�V�"̖M�0������Pw<R��$�V��<`��d�ԼF���i[�ф���b�x	'���~&��H�?C8&������;�:�0���÷�u%��,i}��rN��$�CV�:������zP�;��1���7�B@+ʡ�g۰bq���`R�	����["�j��[+|c���t�>Y�<��e�����6��l?��Qݝ<QF�g�x��^
\8��~�(ki�ŧ��0`��,�(fo+1�eVR����Û�<E-u����<�|^r�z����L�H(����y��^�����0`��f4�M�6G}0G�[�+C����^p���G����:.�m#��/��
-6,�}Qy�����2��#2!����
N�b�R{��	צo�*�:U���P9���_�^��6��7���b5���N<�����cp!��0��O����{�Ǡn����Bu��X\Ab	�&!D���H�թ"P�P߹^ȧ��ڛ�A���$����Vx�@�up����F�V�o�&|�Z¿���$�m�^ّt��&�+�Q��L�8�+��[���&���p|���	��.E�++������6Uu��ިe{e!��[�=yj�����F���� �y�,@]� SRf�gw:w�����������-T��L�aC��v�w¹��?	��߼���P�t�_nN%.����Z��l�[�u���=.BF�nM�ANte����c�	����&�dW &=L:Yz��np�+J�,e�ȹ^	v��	EN�lG�V^�tk0�j�M�^o��㬦I@��k�e�&��x2/%�9L���|��R��;��O$���@�qHѴWP��^���7v��7���ZS��%��Q�
D}�ɒ�~�ݮ�W��{i�k�>�K��j�I�d�́XlxVHYEB    fa00    1b30�V�����ʞ���w�e=n~dZ�Y�Z���I�Ol�6��gx_��h��Yc�A�Q�3��>mi�+��1�X;p��>�g_��g��}���bᮞ~r%$,�$����T$����ް4�d�]��=a���� 7�����R9p�V�-�+�����������Q{䐙0f<r�%��z�a�0Q��w�@�hȷ��H�..��u*:O�'���s��z.�#���uh�z-������iCw� �+9�! �!�t��c&�5��@����k���ݡ^��y����m�E~hO�~���R�#����3�F�i%��"�pT�&��O�QU�
gf�E�_+��37�ҟ�ۛ+�e���t?����M�o����m3r�[�DS<B���U��'8�"M�tD�<�R`(��aqw����hv�e7x���3|rz��4� ez^���*&�i�"0�4�\�3[?4}�@�}q�^)oQD`�Б{b,�\�LM`DԣH(�%� 2��ٺ��21PB5�����f��o6�Q��
'(�@�'Ԩ�i,���	y}o�,��m"NΥCU�����t��hob�O�C�	F�0�����i
�h��v�o����걲i��Vv���,��~�4�������xR���8��o������@pc��L�����w�?��Oz���8̨U���?�����7�$�F��LK�9:I��
�oE���ɒZ��V�HvK���&	���*ܸ�|DQ��(��ؗ�MTV�/��ODmZ�ɐ�?Q��5g? ��1S���b�N�8��mo�7U���� .`!�{��Bթ��$�q�&���jI�+�{~(��n��DWn���%�f��\N��XB|H
��G;LJ�OÕˤ���v�_
��m�f�Wo9d3z��Y��i�E� ������$$�_��<ϙ^O�$uD��8����l�^	*�%Eg�Ly���]�s��S�_B����ZS:S�G��:Y�0͙�H�[� ������X����c$�:<ϳ�BOIG�$���QE�}��zsY����*9����)Q(1d�hA���m�xȮ*����u
��C�N�By:b�
��_6t�g���
D�	y#�^�0ۏ�&63�7K�p�l�?VՆ�p�K������ʦU[����E�3��zN:��s�;� �@y�T�,Q�8+���&�G�)oO�]l��	,L/�m�1����{�0pAR3��^(�>o��hKV{{kҕ���k��9u�H�����(Ӈ=���չ�$�g ����11G��a���I�`���/*\���o7<\%����g�`�?�U�g���R��)�{��%58n|r_�n�&��Eb��_��X/�vr�t���'_�u��k��(؃C$��cuE�PgG����'��?�&<���ٓಫ� �����uEq�w����KeR��kc�1���O�f��;+=�h&�?��o���Ѩ����?S������D��t����/������q&B��@,|�D������;��N�㸐���FNM�����#O�@�濆]q�Ekq*5�/�I���$$�����,��Ո�FOG�� ��2�i��I�	��0�z���\~�8�; �@d���y�:?S!i���߯�%�P�}	Sa�N���#e9���mV�(kW����	���T-Z��[�M3�)��Q8�1��C^�~�����YWc�E|�pIA�yʯx�Z���-F=��U@��m�#����?����C�H�0S�����#m���o�,��;[I`�
<%�-��D+|�ش�S�R�
�k�����T~��U�A�<�x,���AC�l#gӚ�[�.j�D�դ�m��r�;L� �I��*�f���]�y8��:/k�x�´�N�$���,�(�AC����2M
�T�P��
�w��]U���)l��O!��S�ll?
�!*DG�h�����e��0L���!5�Ԋ���J{!�5����V����ۥ�[�N%�I��@����(VSK&�4�C
��\�)N��SY���P:$�1���f���	ɓ��qƬ�#�+I�[�&���J��$O�4~�i`���,Ee�G ��B����(D(���#��O���א+���h��g���i�G�s�s�@*{m	h��B�f_�����'J��VCS7��6�#ɘ�֋I���ÊQ����6U�??_� VC&ަQ�޶�r�N�?"DN��h����:?n��a
g�f�)3ݳFV��mR*õ�a�8�}�.�B��}��S�M0�j��({��}8�#:X�7&�d�ʵz+NQ\��\�����U�����˒5��FU��xW��t�
������0]|s�+ǻL�k5i��Q�α���|i�n�lѪ����U��TQ��6�׃�Hg�k��8�*v�#�8^�6����߻�� ��ȡٷ%ڿ��K�3b�-�=����xk���]|!ן��,�d{�;��7 `:H��7f"WX��
��A��Br�;R�v?v/?lI�d�j�nn��d$~q�$ĥ����7�)1�WB�s��8EO��-�_��SY�?ʜp9\��Ϧ�۪�՟�M�������5�j�+���KPK��V$\}Z�-qo��Җ�Vȍ�n=�4d�'�G�:a��/ճ�D˪��.�7��Y�oI�j+@a�\QI�7ȟceN�,N�G����x�P[㭰 �X�m~��̱����P��D-�;�S���1�S��"���U�]u��H��B?�WD�Ƕ�D��Jpw� ��3#(c�'O��-��� ��ډ��47,�=�&W�ؽr���H�o�C2���M��{Q���Y�]��~a�* t�|������<D��5��#n�琢NSa�8�k�jf�J@�wb��=^`�Y����sxf9��b�ݥ���6M�~��&�(r�+����uti��*~�\ۃ��8C�*��/�BUR�Bp�#ݒ�#���*�B>h�Eޢ�l7�B���E�e������'Jg?��~�G�k��g�f�yh�w7�Z���nC1���H����m�>�پ�Ϙؖ�}�{9�5���FT6��Gc���vC
m6~9����B�gJp��2p�j�����=}��~���2�GH�`>M�8���9�]�%�-��K��VlL�ry��:�ث��3���B�� ��e+�Oj�zd��� ,�lr[W���PV�RYu�����~�3���$s�Rt�hp��>i�#lr�=d6r2����{���)5z���ɧ�84�Ł��N���b.m��e���N�:^��k(����)�W8��)����4�Cd�,�>��~Y����z���J�m����N�&��L�Ji_�5���9�}U,ܖ�Y��h:�(�RYh<|e-F$r�v�i�2����5��Mб�?��[oc:����ԅfΒ���aV����� �پ��os[�MI(�>��%.7%C����%�'7)��(�ڟ�k�N�5O��q�,�wOٛ�yVw����TN嘾�4)CT�6�8	b�֠{�T3�9�y)vm�Z�j`d�J:/ÕVU�E0�$�evlD�TN���7~]V�$��F�BQ�;l��)��Ȣ�F'^^(W(쑾97�T�$6��F~�Y.G.�75�a�2�K�4)kɥי<	6c��b�:HYr����^��eD2Z �%�.��Jj ��>h�p�4Ga��!��6��vn̈́�$i�9��0"يh�׶��i��Z�1�Q]�_�j1\?*�~��V��˘�GJ�VC�B d�ͼ��=ҊЍx�x�>�<�t����6O�*DE6a8�o�����Qs4��h��%�¹h��<����30�P���ּ�����CP���.��#e��&P��/���&��de���Idr�uLdG�	�ø�.� n�6��3���3�WQ��{�b���7EFi�^�IWe���,��l��֐�Nm�5w�?@�>υ[��[L	�n�I{��T@�"�F!s�pش&�9H����3��:� �0�JO�a%߇��`3��P��9�q�]��GV��.�[�e[�_���@�Y8ȸ�����g�F�d��6�����t��CryD��ƈK��X������p@�A挼[���
y�V��>\���B�,�f���=79�Fƃ!�si�Q~�c	,�y��խcB�f�e*3�|8~��I4�q���S�A� S 7�ה�#~C��S��v�Iy���j��Db[���xh�O�r%��HZ�n����=dA�#�(�U��3;d"�܋��2�^=k�
��s��MLQ"�OW'w�$�����oO0��'���{���t!���q\.d4������z���n��k-��������u�Y���	w��jB�a37POv9�<������� m;�M14U�R�7���f��2ڸ�e\O�e���5j  mB�X��lu^	SC��C!#�</��;��;h e��S�ܦ�C.���,��T�?�ǋ�v*�m���d�R�tE9�6�����(N�h��g��[P���ɘ/@y������*gG���	}?$���Y�EM�+�g F�Q8��Vn��'�7����觐N"���� ���O	�>K�ܡȢ/V|�����U��&��en;�%I��]`%�G(�;,�e'/�1$.�ԉm���\I�P5��ú����u�y˥�du��H�?j���� y�׽rx��&�$�����;�$<�S�L�y&��
�����fW�Ȓ��5�Lp�3��Y��y�86�5��=�t
�y�
��XO�T�
�b�(�q*k!�k��mW�q<�:��^ͨ���2���D;i�786���;O�u�[�&�r�n"��0�T �#@O�S���(,��7
%n\CU���(�	�N}5Z�қo���FϞC�����1�
 �yI���*.�&�Ms�N�J��i��?�Z"�,ʊ�{J���^n$H�a�r���7�51~�؋���V^����%�x:�+v�V�� $���yTM������ ��'4��ms@��h�X�z�~@��
�O�m)Y�˟�m �0:n@�M��:3N.��H�O�W �����u�?��w�:�����weKR��m/*�7��RR�S�Q- �_����ݚ�V=��S3R�N��� �,��������"�q�f#m��O�k��VҰ��HZ�-�m�k3S����"���bv�C���4�	Ls�P޿�*��=7>g���V��{��i��Ym0�)�F����5H9S������4����f�3��-x�}��FDF���<��S�*�k
�$�=�l�@�a�������W�'須B
�s���!��$�Y���!�׏���yDL���]E����30�Av?O�g�����JA�E���=7$R������^��PTگ�I��Q��;���Gx��nP�SS;an��\yl
�1��{HL����g�g=�t�}x�gl�d2������6q����*k��tan2S�f:���:����1����v����c���q�8��%C3�q��� ����a"��1���EW%|W�~��o���g��%*���܎%4����-��2��j�!Ua�D\c�$ax�J]�Y����w��注DhG���܊3k� ���=�ǷB�I��B����tMQ�ew�,k��ɘ��RvZ�\�)�����l2��	��(Ҙ� �<Cށ��'3��H̐gVVo�-KT^����1H���:+?"��6�D�'{�6��,�S P*��U��pL�r�X)^z@dGՅ�Z��,0�RZ1l��=Z�S=��衊���j���"�3�\)n��B־Yб���:��m���U�H�k�
Dk@�:�%ʍ���5�[�0R~�%���:�(�a'����V� k�>z�{-_���d6�%&o)jxC��5����}��L�P��C>e4Y��t�(Sm��p�)3NB���a�������c����\�!������ԉ$����:S��%3޻�M/pM���T��#я�E�#�U5r��i?�3���_�7u�նQ)V̽�'��6�@���HS�H��_��2��d�О��-b�����?Vk@loZ����Q�(١E�TTIo�����{������4и�<��5ֆS��Ɣq���6㳐\��<߻A�'�8��Y�y���i���8������
�O#�q��V�e$��C�T*b�'���C݉'�&t���}b �Ӭ��c�b7�s���{m8�<�(�	Cd1ϛW�SI�g��a�y���>}7>~ȁ���]+�-�iu�N��mI���f5
�n�sJ�S�lD��Ѥ �����NK���/�.���*�B����?d0�^������)ίM�@��E�v������I�0��Z�����
��a{��V�a�*p�	�C�&�u��ͽ�<ꗽ�{[���g$�F�e��\����U��cţ�}_wC2�C>`�j���
Ę_h �Β�=�����Y�_i����Ҧ.t��]Y}u!c�0������*W��X#�7O�v�5�ӿ�]^rS���B��RzPV��Ŗ���ל���`�X4�Uz���t�	�΋F6�W|�gm؃F���҉l�r��'P���Ҍzgǰ�3��#=��|:ӠǏqj}m� 7DA��g:���4�5�!ӗ\�;�]�|W��G�!<n�X��_H
0�0��v�2��HcQ�(�(G���;��C��!��׆y���K�$мӠ�r�����
����Ne�6R@�,�<��ް�36Z�͓
�!8����c�O�U�r�)!#�/N+� tL]�8�Ǉ$���2����(�tl7.U�,�5�U�JXlxVHYEB    fa00    1950����:��f!�5{��[���/����w5�0��K"�/�I���R,cI�K ����
�.cE�CO��� ��X�����B�{����XL�$`k�ZCE��a�]h3T�ۅp&y��'К�؊��lD��z�4�Y��aۍ+Z�i�0v����-���i�����:ܖd��LR�"8�>{q3�w�P�xS��sk�눀Q���E�{����p� �q*�xK=�t �c'�.�n�K�����y_]�WёKBm>�/��s:"��C�.�����6HƩ ��=�d���Gk	�Y�Z�S:�G��S10y �J����ד +�5t�a�+U�״��b�מ-��X�
�x_�uW@�� 2�9��L/����T��&p�\���<*��VI��j�T؋��Ӄ��A�?dzd���mt` ��m�N��Q�6G�I������׸�hX���:��P,�l�f����k���9����BGիr-+���2��0eu�֛�0�f���
��d۶�Qԕ
aw��UDn�F�a�����e��i�|�	�S�G�3IB�
cbNa��n1^uos#��h�.}�^�z�1T5�p����h~l�AB$��讎'�;��1\k���7^A	�%o�^���^���}�j	;���q�9�R^#d~���^S� ��.���G�lLh�"ޯ5yu���ֻ�Jf��c��Ȱ�7�({�&�E�7�uOJu�n�����Ӕ�S~�����e�4�=�X�{����B�&R��,��5�Ǚw�82_�B���Ӹ��-�ߵKl������p4�m�]�=O���P5)V���g��@!��w�`�BIaJ~����[|U�S�-�<�j���A�z�hr���ݫ���2�K�9�SJS S��oNi�AD��P%u9��_k)R�d$�6�-j'� f&L<�� -{���\�Y��X�"*��7`&�S4�/%��u�%Q� �P|�8��*D�&w�����ί�B�*�+���!��*z:�������To%6pW��wޓ-Go��y��$��!azqݰ4��������c$u&9�5�.<�]���T�i��:h�M���[,��	v���_|�^js�"�Z�$߯��)qÑF�����/ ����ç�j�rM��(c6�l�����(L��������x��U?��s�g��^��捄b�;Ѫ	�^4��qQ:XX/
�{�ѠU���!Q�U���@��6�BPB���=J\N\e�p%U���!*�ՙ��C�Z,6�ڮ#2ńKB��ڪ[x����ݯ��h�O�`-H1���yX-�x��5�Y����J�)̖�y��z��JB���M
��D8�����*��^�8�o	��u<|��O��H��ꪒ:��27�#;�>!g$��*<_�))��a:.�ڲ٧Qm�r��K��q5b���a�^��U��x��lM��L�K�ā�b��܇��ёb���RH��W1����'�5Z�L�5N����-�.�,�z ���xM&���Z���q��<�<Fՠ�c�ة���/TH���������D)�J�dBv<J�\>���#���%����[+�>lZ]zH"/�r�W���	��+	���|�cw$�Z%���zdǉ��|�]=�f�3�<��l��z�_���k/����9�j
C�,���,�S���i憡��ǹ̿��?Ssba��� �y�R�u��u>���W�^{�>0��,��b�����4= �< 2�}_�Ղ��2� ��Ef�R�:\��V~�\Dc%[gT�Ğ�:Y�4e���qvf��ì�}J��T�Xmu>�e���H�jT����fˮ�@{�w�~�'�����ҋC`�-�<���k
�\�>IJ#@�v�!��ؑ�t��>���X=�)p��e^��o\�����_hn�h�� i�q�\���E�_��v,0������cH����>�m �\���c^C�i��J�b�HRX�˱_��3�n%�-t��y����*pi�9��	��gT����VL�e�R!ͪQh��ٴ�WK��W�k��:PA7$0燌���;��S������=��D�BM�B�ƹY���H��؈��$Z��E�S�O��3t�B��}��h���C/��B�:J�N��z���3c�� �YG�W'g��:�+�I�	/�Љqu�\O���)���%n#�S��䴬��e�(E�j?-�?���;�lаnu �7R��9�Hc��3bI�O4�\�ä�nQABQ�M7T@�i�G�Y�K��[�>�=T�B�M鮿57����u����Udѣ���xf��f������+�=oj���,7J��Ǯ��%���r����"Rz����?]D4kE�F��6���ki-��:�uu.�#qf���� �ͤԱ�)�g��~��}H�D;<����x�����4ĝ9C<<�Or�I_8�h�JE�b��L['��ی4ד�;�WO_n�ز �Uހd��c�ȩFx��8�N��G.��|�������P؞B<�1���K:i�iUR����r�2h��K5�|��-��WD��< ^˦��v����fb�<� ��v@�Lf�a%C*$�L��<��-Q��,XX~�;�+BP>�T��_��7~k����F
gi�RX�=�5wYk]'t��,n&�Bb��׵�GܟB�"5�"H��Y"<|�~��a"��P�uF��L����r��S�Rf��d+�8�;��Bpf����|� �,��If�G ��p)����x�Eh�0ðqXcΗ�ķ�&g4L^O�5UB�ڤ*�	u�h��b�o\y�lߓ������`�-!��3H6�h/�q�t�R;��]	���b���>�c�.��n'dǉ�7��X�/���R���\�[�>=3W��:��r[m�BaPx��m�}A�:��(G;�q���]� TJO���W���6뗆��ѥ�D(H-���?QY=0(�{b��[�w 4����@�T�i�"7Qb,�i`��G(�I�Ki�dj� |��Y��,SF�Ŋ��/�y�Nīe �CΎj!�whB8�Mޓ��½��fV �"��}Tص� ����4&���z�6U��=��Qc]��8�t.x�65�~���jc\����Ң�!��t!�9(�pK(�:4l/� d�L� �l�N~T�p*��D��M'sHq�Q��h̴�ևsy]�A�i;�u����n9"��1�z�̥"��C����Aԇ�g&��1�3m�����5q����,�}c_�����R�c�C<�z����������c�i������MRB���"�^��y*NL �Y�w� �坩���H-��,
{�������aF{K�o���3H疴vǊv�78�&�۹��?�"����H��"�=�*������;�]���9��@ztu�@-����R�k��L��J��������ӟ�i�i�V��{lk����쳸��~*�Q���4�Pmn�eR}�!ij���7��R�SBe�"��8��V]��iz�=�lv����+k�2e竩ltRX��P�E�W��M,�I��� j���o���uϰ1��Jw�O��':��v<Fg�~b����%��7�%���m�xM�����ٍ��?�ş&�������U]��_����?x(�9�P%��O�F"��w��Kz�_�?��N��_�I���n��t���,��̓&\�7W8TCsP�2�B��y��N�W���@f(��=yt��� ��u$��y�Nd�����*��eW�q XGg��`���%E������i5��a�텊v]����W�I�V�k�/޽ Tص�3�zr�s[w�bkɨ����&�|���:��䒧\����g��i�\p|؜�tK��su��Y���)K/���R�i	��R���:�8�����u���<���۫�jOM^���n�mH.��
_��.��$A���hx#�ӵ�z�]�:���P�_]�RBk���3lȽ�ɋ�C@����r�� ��3wh�~��E��q��9�E�{̷Pd6�����	{�)��M�_&��!�J��8�b�'�ƣ�D�0�s�~
�B@ND���r,�/��t�R�&�S����@�L巵2�sZZ�fi�wk�AI̝o<'`0�n�-L������%'�c���Z-����>$U�RK������[����A�a�x�!p�8�#�Ǭa�������#��%Y�_�V@�M��P���V��ᖮ<���(�n!��ȴ��Եw��?a��p��:W,n&�sb	c��N��Y�Q���N����;�n�H�M�Kh��p��x}���%Ř��w�as��)Y�pga�%k����-h��uNYDXQ,i�鲧q�q�m�����|�#�)�I���ڃ�G+�L�Z�u
Rox���*q��G"������r�F��a��\�$i��善"�g��< 6Ło�F�(IgC����������v�T����ț���N����X�:3�Y�5�[�^K�!��k�Z]u�ع�m�Ǌ?���
���OE.�a�!�Y��"I�<��1�F�,1`���'8=�/�g�oNNiK<j���yB��~2C,�@wt���n`��qE��U΂%q{|�[1�zM�qGѕ&���i]�rp,��&�>����4�;��#sHFy`3̈�!�C(�0����F�ʫ^�R�A�*eJ~����F�%0����ƞ���ؖ):>hJ4���G�y��5�7�t�j������&OL\��7����bW]��S�9���\�yi�@��gJV��J��c]��8T/P��|D�ْ���Kz���,���v�=k:���"v�{l��������4s��u$F3���X�ק=�~ۊq�h�٠^��Ϊ���s�����E���/`R�Q�	��̧Y	����Y���nJ�q��S=��c3�F��C���0F�����|�IUN�!$���G�cz�`���+퀜`���t|C9it7�/c)v����ya��yV��{N����ɜA��U5��H�⫎��$�M�&�&R�<�mɿ2,�|�xy�u�Aq/�-/:����O��c�_����T��c7�M�<$��qfE��s�o�������k��*��oZ�Zܢ��{7:��{�8ʂR^b�2�ݳ�M�;���C���g�G�M�hiC��Z��jI^2��2��i0�Sl�䳐eF��T�/�C��=텐���rF�	��u��;=I%�~j�%��~!�ge� *�0��9���-_��}v��
;��9��V��.Oa�І�f��@�6���ƀ.�r�
��j��K�^r?�*� f9�vv!�(�F���0,h @�lo_K	@�����2'AZ	E�{4e��<�S5/t|�3��{0��4˼���ppR��,]!����)���gf�DW��n�K��~�z�S#�f7-������+�3�F�l�{�;F�M��g�f����p����"�D�T���0۰�!G�J�n��""�.X�\U,7�e�sG�}�|c�z\��"�M�ʑ��fH�GS ��Ҕ���f������� +�nr\�N��+GXQף��A�F O��&�Q�l�ڒt��vW�c�ҝ�\�G�a��9�J$�_�������DK�7�O��T��'�Bo B�V�ӛ�/q莀�]��yZ����َg5�W�K{5�zv+�g��������H�:��5�@�W/�����@vsF�i ]����,Յ�t��0�� L?�G��ռ�]6`��oL�i:���0�Nn2�G�Evs��I�gʂ������0���;ժ��el�	��3}�v��w��f�yPOam6=�lN#�j�Ԝ�0M�b���Q �f�G��:B�䩁4�X��<!�<f��H!�̍^V�l�P�}�%i�&	.��{W�"�(�6�G)1�o`͝����Y/����̶ni� ���Fb�'�i0�4�å��
�+� NH#$��/�!���u���}ޔ���u�bE�昭��*�rwx�&·�d?K ycqI���ڮ�g���L��bՔ�i��H"-_m�8	tDΐ��p.h(��dg�qU�f����3')�><��e��RjB�%��O�U8��u>d��Ok�	���@' ��
ǲ���dzh�f���vw�.n��N���V(TEL{�����n�fF�Nm���Z�ǡ��#{��CO�5<pO��s�xY�0���	@A����_4����}4��"�i���Q��t弑$�2߶i�0��Ҹ�d?�M�1l�4�����9<��������(Z¡�VtE��h�IWi�XlxVHYEB    4f3c     d50
=�Er뿊�k���H3@N�݇Px��c�a�
����Wu��
�̌�� /���%_�4
/)R��j��%�Z_��>Nw�׊��{d�`d�S���F��К�Öa)����
N6��@� ��19U��=z���eѡe�zVL�RȲ����%jo��Վǀ߉
�΄hmi�7/���<�ֽh���"@��r�/�v EU��R_��"�i#z�57�A��/��"Ew�r?u����M�ˮ�EP�Yu�'u�I�����b��2G���&󲎖΢#�� �Z0?�̲&��FF���}�|�
V����sƵD"A��ȸ�,x�d��	�����b����p[2����l؄l���Ff&���Q�Y�2'Y6���W@��y?�e�󢯪ݕcr��0s��B��V�/�s ��<xv�|�m;�|k�df��~q'{xۇ�gs}�q �9eW���/q3(�iB"��ar#a�Z�����7Os�j�v�00t��A���:���ɉ�b���iv:F���P���/=3K�a���,|��Ǡ��ơ����T��8�2ݕ-x⢕A�&��6K��߂q���=pHH�ݮ�dBK>���G�c�]����k�.ag�Ա5Hn�������é��@��8��n�p���N�EQ���ߺ:��OJٜ�]Gw/�m�������~KI6Kf]L`��yc)).sm�c�]�Ҝ�ͥ�{�"B���1Q2jὟ�[�k�J���W�/�j"��Z�׵��V{G�UVULh�A����Ovj0��2$���M�� ���7���3�
�V�d#3�D��F��s�~ڰ�7�M��699G�ǚZk!Q�uʯ� �4�	ɰ�78�9���k�>Ւ#!� 8�B�S���1N}M~�)�|!y�2���.���s`l&T�E�NF��dVi��gh$2�p�Ca�B�* ��E#��(�PAP3��~s����1�=�ϻN)��c������L����C��n�r�$CY�V( ��Ź���7bB=�M��Z���Kd��% ��������@8#�}f����`�1`�� 	�j*G	��_�r�3�h5iyh�f��Y{i-���s�g �q6�.�ո������w,S�Xr�H���`��3c�o���1���a����d���������ܢ�j��WJޑv5�˼��|DkB��~���>p��3�0 x�gB28Y���<�	�
7���|�d����6	�h�F1�F������,��G�#�V��fф��"H�Z�{�ǖ�◧y��$Q"��WGs���dB�d*[(%��NIʔ�5�Ī�����x=X""��bv&>�-�i�X�;���>��/��4*>qZ��#FC�Q :2Ԛ"��T�?t�j|!��uEOێ�kx;=��F�c��a�V�CJ�S��[��5�D���b#����24�*�?�� |�����<���I" ��`�z�-bUL%��/E�^<Q��;Q�aC����-�ꃸ�D~��g�z�8���gbG<��X�B�<�a\S�C��w�K.�Q�֭�n�juu�R��J����/����}%g�S��[p��x9&�U�~k�rs`��^��>نH�L GU���<m$݊���XkX���j��VGVH��@�p�	��m0R����rΌ�e��IF�͋�x�ƙr���^9�赉��W����^�3%�m�
-��w����G�g���ׁ��EE�Yѵb�d��!����qt¶�@[�\�M�3ߔF{����������/D�Y�sU�o��]`4�e��G�Qȡ�ehY��ʹ�p}�3�6�0|�a��WT#���Q�\~���)�Q��ld�(M~G�V!?���^�>�	�+% ��K����^t�B���1�Sڗ _�lCJ�V�Qa�G�q�h��LNu�Nf��a$Z��/J��b��-�w7����$�?��f;#��-�KG?�qO�sB6?D�nM,clKvL���?�:eM�rW�\�mk��<v��m��s�]ʷ1�6�%n�j���	LlIG��b@�Kc��7}��*��3�ۃ:�q#�r���ɶ���f�F�ʄ7I��~v��`�v���g��=�;^�H�`mg+�40��'�6�_:6����T�
']�sL��i�ӎm�&��p�!���qZ�R�K[Ay���3@��Ï-aD>�j�u�R�2���QF��.TxD:�:.X7�� ��<ٟ1��ش���>a�;ㅊ��������[p-�"��pH[e+J\��h�(Z���ԘD_V�BGW%���
�_��vR0�.S"N���E��?�1���
;��5�������Ƶ��U1&}:F�̬Ŏ��S�V��e��H�3�7���l߲���@�%U��Ӥ��O���-�6�`��w�<�_3q�sm���u>�|Ms�s%ݱJpyWp�&�	q�,���Uv�������<�K thPɛ�@���д�U�lR���٬�ݻ^���8���/�G��sr)h[�c���"���v��?N��G,�1���9 ����1���o��^��5��;���=T0�qRa���Ѭ���],�9���$+�g���EM/A6C�q��ᇥvjHѽ˷s�ީ��K�khU7R05+�5��lqsP��Ӕ�v�
́.�e�٤rv�k��5��ߢs
P�A>@��,l�����t;7^��n�\J�����5�]�w9������:�~�Vm�s^4���`.d۩��)�E��)X�/��#,����Z������ԭ���I>c�n���R�P�C�@��gH��?M�l�#~�$�Ʀ����Rr?�v�V��2o����x+D_ Ԟ���<���T��\���8�2
�U�������2�^�F���	.����k�\O�K�{��7�q�U|gf{w#AZWW��d�J Λ���]���"oZZ�߮[�����l���&_!|�i{��W�	6F���}�S�&(��u�Ho���Y"`A�OT������c��y���k�����Pl�,N���j������
��l������k���F�1���wq�,�o�yxBN�u��*�ܣ1[E� �V@�Y��~D���8,B�23�/��|dge�����lt��/"�ܯ�dkR�Bh�L���el�x���v�/2@e?_0���W�{��ғ�s������0Soûnn�8�(��ԉ�8+��;�&s�5��k_���U(%���s��`��yN@���)ݫNޝcAX�f;b�ҥ;�c'~&;��c߂����m;�a������M�V!�+li�O�O��^�b������t6��9��x������tF$\��o�ZEǾN����u"9�Ǎ�܇�Qf1�{�tëx�Z��$�㈸�¿ɑ�7�����Õ��It�t��!]��Y�