XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2��bX����0=�Gu���#k�4�&�h!�N<��\��_���ж��~�8�bQ�o���l�0���O���309<A��3*EJ����XS�C��5��8�4Ћ�m�e�G���T���х�א x�E��o )�;���M�e��~�(|X��+N�3���S<.HX�9��@uI��M���HNYy*��zQL�*؜;��S�NMs ��q��0�K?�������UN�5"x^"�MI68�rY<H�3�]�V2�&��Q�o^�d' 
J�����JT$�6"��h�3��t(�G�x��w�Ս�3Z-V?�J �6D�>}ߡF�#M�:(�B]�+?˘7$�j)O(���x5�y��C\��p�T��4:�g����c���b���t`�{ȇl��Pn#U�N+0e	!��LB� �0L���3!w�I�j�Sp=k¤�#���|`�$`_�ٰ���{��禹���fϳY�J@���s�{�N=�|�U�9���迵[{=i�B��n��^�8 ����J����3��P���:��~s�C���Z�Rq.�B+�Jߛֆ1��n�+��B�&�1yG�پs�"��X����B�#�I��X�q�hllK�;�ɽWճ��3�2f������W��6U�d�FP���Z�_������:Z|�
��~2�g �����X�}���y��=l(�ߘw8!�g�� �݆��u���v�D�M�_p?�w֥�ں_~`�3\E�!���[�&�BW���XlxVHYEB    9732    14d0'����#�Ԙ��p�)[#+���f~�w��E�����A�R����FU��1v�	��D]��ao#��Z�+U����~5V}�R�e�a����UD��ܺÉ�>�F���6�J6�v��>�:�c���N붖��dޞ����H��u�43U��|%�E(���h�Q��͆� �rIc��ت�:�z+D��4����S�0���g\-.aj���dc�1J��t�hREⓦ�a��-��6S��T?���+�"8��r�/�k��z�g�Pr��n�ʜQ��	xO�d#��-�򊔟�,X0.(6��������1���׹0*hy*�8���,sh���'2*��{$ǀ`��І��t��F�/�rW��bb�T*��N�t'�����8�qa��}$vJ|?��� ��PB�BZ2��DE�*�e��(b-�U���G�	-�X��Q��c2�lƩ�t�h7��q�?}�vұz�Tg̹�t����F@O�!�"t3��T�^Cc���`]9eV�?��W���#5��*�,Ρ�3/3s2�`�;YPx�W�{C��S�� =?�Ig��_��ǯ�r��e�f����4���z ��B�C�ڜls�3q>�R�-ɯ~��dB�@j�[�!w�Z�d6��� �\jo5���7�l �Z�2ݑ:7_�"�Ҥ]���(�F���	:i���/��g�MH2dw4��:�<8H��j�p�;�]�Z�ۚ�H��������v��J@��8x,^��y�dħZL�!`�6��=��raSB@M�x^Ecՠ�O����� �����Jkpi\E��ĕ��^��|�<�#��/cC%_��-@k�>�ӟ�$[�q!��PG��GZLM1v���R�0ǐ?	�ѓv�2`'�Kѣ�2ё�Y��sx�������+xr��M.-���-�b��X*��z� ����P�a7��e��t}�W�;Kf(���@{G��o��w�� C�JL���ފ?�7� ��~���Ϳ9AL��i8�0�:�o!�u BH]c'���v�䫦�Q�,cXwz&"��X����
�����`�#;��g!���j}h�B�:�F���e�����*b춍ԗW咺���⫝ ��� qÉϹ�Gʕ�o���D����ޏ�dJxU�鑰ωo|r�ҹ1	^ MN3)�|+�֕^q�t�_���m�6����_xr��ť��^Ӌr{�2B*_��T4��.��Q���_��Q�ICaT��.�>χ����
u.���	�$ �D^sO��J=��N4���ZF��a[�$�*Xwh�ܣJt��� ��c��S��f=X�b��Q\AwM�9|p��?	C�v�a^V��u��xVY�L�Lk?W��#hf�\�Ϊ��+�@B`h���G'��h�I��,���D����r���m~[�#^0���Q��$G�f'�Fe��F\�Z��ؙLX���k�-���K�����Ձ*N�0��dvM_���v��n�<_���[��O�js	M���������П��b�Te�[GX�C��O9h�����R���r�K�\�TErnQl�m�	(/q���_[�:�堙Xʆ��֤� �I%9;
r��������\+=\�n��ךH)�sj�qo�+7�HfV./pƿ�t�cbx�{ܝ��bW��?�V���n��W�\�<���m7�>��x.�.az���jS�K��ik\�ա�E�,z�U(2@LCG����t;J��;��x9w��+`ǽ���6dٱ���vW1DQŠ|�c���KٴA�׉���ȁ�(��l�g�`1��TrlÊ�3��
/�^�H�p��%Dn��_���g�&� g2w�|Yg��8qo�_ҕ�:�+��j�LQ�[`y���H��Ʊ���8qe��Ȟoɒ�����'�1C�=?��؛_�B}S�3r�~��;~��f��Ѻ�b.ADqq7/�z�3q�a���RO��Ъϛ�ư�?�0^y�m����%pO�{H���T�Q���b/ƍZ,��S;��1�z*w����4�E�����~ٹAfw�9@���Fڸ]��i��zD{��~+>o��ܲ6�O��7.�>�����
���y���x����z&A�"Ygh xMF��!޿gʓ`jr�[WD�PfwD��Xa��.�f��WA���-�n�Z�^�	�Xw�,R�R�D^�ˍ�@m�2D3?�5�hGM�R0~Xb��"��~�K�4.�cbD�B���� �f����o�:�H:�0��	����*��Ƈ� ��E�f��eJ�����so�EYg�ʋe��Z�R�md�h�/�-)Aŋ*&ߩ��X�Di*�X*�2��=�Zک�)�fQ��ܕ�W��fg�2���A~*0������v��.�/�R��M㈊�Lo �O��5���D�� �٤x*:���)������]�"�%��*w+3
��d|���ؿ�{B�+Y ;��������uO����ų�唄��NUB4Ф�:������r脅* `��Zl�&�t��zu2�;��X�3n&��@/	A�mF�/�{Ø�'N},g�ӝX.AT��3	��sJ*%�|�����<��
Յ���;�2P sP�:	Ծ^ #�Γ`�y�sr[�}Y��Q��*�q3�Д�5O��H���_z�a���$,l�4%Tj:`O�^1#�?"��ΖS�&�@?�X�� Vo�D�b7[m�4�<3fQ���.T���i�꧂b�Šc�����QP�;���BYCR<M�Z�A-j�ӫGa'7v��QMo�Q�|�EL&�*.����Մ9��t�;Z�f���B��8��z�S�GL����ya/޻T[�a`z�]NB��
Έ�1���pd�e���S�mF��!>Y5a����8������m�g.&�oP����%�zj��T��[������kݼ����SJV>R�澭��#|ZL(e���0�����ٸ􋿴�$�}zc����'i2�6�gkHBfi��TA�)4��@+���k����6#��l�@���zf8-�I=t���3v�D?�Ac\���4�������1�۝�H�R_~��mO@��+9�<�6��)�R6�܆�:ѐ!?��LZ`�W� =O�n�&����T�A��`�w��[�4sȎ�_'�O�Ⱥ�|}b�yտg��;mlx���K&Z]�B��F���q�&��l:�v�n�{�x��-��\�7s� W�8�#�<��l���v�±�*�VMf%rX�b��S�46^1��LpOtD<6�`x*�Q� �`h5�⸮���͑t$�SS\����H�fg⟂e��Kw~�=k�f3j��@��G+~P����'vG�W��Yy���mp ��X��4ɸ�1��sarE��qr�#�	E`�ݳ�{�{3��[�^�X�՗�v*�l �3�yn"㦯X�6J�gv���0�]���i�Y�ܣ<�������ܿ�q'\�� M�O��P�Fa����v`���HDC�2�鮥L�L���hMS��f�
! _�֞)����ֱ�X����1�̯{�{<
<n�*Y#<@x�pk��*�FI��8~L��'�c�Ӟg��p��3vRs��+:�n�L\�����"��Ԇ�i���Iv���a3F�@uؒ%��垱0a�����yQѬh�;Wc$C��'��Ⴅ�6��jmpmV���|��v	�5�=����h���ɡ fHw+	�J@�Nٚf��~)c���(��s(����N&^b/m�黰Y��|�þ<H�����,H���� I;�:rI���|��o�J�t?��)6�����a���	)�~)����9,��k��Ϣ���(�Ҝ�3�����َ�"2U�K�&��[�vr+�#��(7l5�H��� ���4Gv���"Ѹ;Eņ�gևx���h����4�bv�xQ��Pql���sG��ȱe����y�[�� �5}�����������<�Y��;�� ���{G��PAT��Om��!6|"A�i@�AK<><�p�K!},��V�V.Tzb[�k~pnU8��g����G��K��	Jo洂x��N�[�S^:RN{��Ԩ
a�a¯�2���A�g-���I�?��G�5L�����lٮu�)�v9qD`D��0�dp��<���I�TE���)�s��6�9�=T���; �Hݿ��̦m
1����K�5~KX�6)�x�n�h���yŤ��7�$�u�1e^a�%"�o	f�	��@�=�\��q��
ٰ�֚�$��e�L煓�:���� �IP��	f�ں{��h������d�Ӕ� .���q>�g����:�Q�.�6*M"e ����d��L=ј�6��1���Ğ�ɦ"��, �m���E�⟐
��As-���3]�NG��h��zXpnSz[}ZU��k�Y^ʄ�-�il�;a�Pv8[F�~�����z�y���e�f�!^�>���a����A�Ї0L�N�~tZ��n����W��O�NK�!y��z��{����qu��~]�w�Y��>|�k�F�p���͸>ħ�'.����X�):�<TI	Q?�u����qp�H.޷yv3����-Ԁ�cJ?�j26�v�t0i��t�����	�է��s-�V��^c4�m�$�m��a����%��r�&i-�+�)��Csȋ5(ݛ��qϠ5Iv+�L��ڱy`��Ź�=u8�M`��3V���{g�Tv��\�zhk�8�N�E�x�;{P��1�A["흞�8Q���3���Jǟ7�_V�����w�L5m�h�J������b�RݒՀ�h����"3,3����CS�#�� E��N�)C�"͟<2������=��x�!�#`�IL��ZMx�5�ӊ�ע��6�#ȑ�A�z�FA�� ;�ٌ��-��ݨR_&�u��#+!�`5�7s8�~�u�<�Vt�\�MřV�����^�a�W�2f%�o�
�%O��O��"�K��8����,� [�m,5�r�c��D�aT�͞��@�YTcb���!�N(�*B D7���I��o"25�<Ԥ���wJ#{��\oP@x#�^D;�w<c+��z�."d���:߂��mME��}+r0Y�;�}:��8٣ڰ���6=!tǓ��S��f���Pb���v{�NC�u��)9�01��N����|��`jڳN� ߛj�k�G��_$N�*w[T�4n�nܠη��K�H| �`�"����&a�9�h n��ԋ?�/IQ]�����
�0MUS�gx�]#�2nuw^�V�ByY440