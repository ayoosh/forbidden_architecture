XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t�V�8�?�oY�0��	���u�+��m�6���m��7ͻq1:P �`����8�f'Z߇=�������?��s���W�c�J���44y���q�L��_%����6�{��W֠>8l�[,Ԍ��������6�\��u=e��B��=���ӎ ����+�`7��iM/����,T}]���q�n��̡=��+/�����c~'@��Ӛ����e2������&v���oط��=km_�����!i������&w`!��M��{;d�?��O}�����j}چ>�S���������sG>4��>#�s�j��N��]p4��+��9��NB�|�f�x~o�������#�n�^"�wHrq���}�+��8������!�4��h�+T�G�1�.��^DjC�!uK$~���.��b�9�]�O��vH[�K����+%�����e\�4H0��t���C�_���c-�O��9y�ÏO��	��qQU	���@|yt/���s��S����5Nᒼ�ݽT��'�P�x�h��Q$�򴏸n� Xa��B���z~��O�`�p�����ЌBD?O�a!�W�o}ܽ��vH��F����I����q簮O"���}�:yǅ���,��1��I�{�!
��Y���
��1 H���Y���&���Eq ��q�*�;��g�D���bE�����kOTF��	d'�MV���8���^��*��06�&	� �x�u��s?��0&|l��<����>��=XlxVHYEB    33d0     ca0����q���~C��l6�*?v�X�G�Q�H:�B�F���f���?�L#*B5�KJT����h��XT$� YF'Ԉ��L�E�K)��Že�C��Z���jc��z�QO�����*�aRwm�9'�\��C�X+�/X���/��K_LH���\'g���E�
���$א��z������Bk(��2��V+z�T h3&;�5O�?/�Ӏ�_�Hh��f*v��M+��@�S�󇿢��m��	3��A��N�gl�-��sϬR ��͘���!hJ�l�~�kv�߾��ax�u�!���	p����<b���ˇ�xI+$H_Yē��G2��7iTC�Fm��N�'�o�@潖�ȭ>�Lԁ�M�J�Q�+����h�<��ʆ*۽u��K������ ��h��[z��\�՜�a�^>��Az�j�?���.<ͮ���<��w#�6��x�FP �.u��d��N^�M�0nρ�������xM*ҿR�UW��QRܶ0����
������#�3�Q�XG	H�`���]s��p��푹�9��#X�BǤ3"����/BK�i�����.i���},��~��<���(nv��<lƸ�T�ʗ����(I{f7�-�KTѺ�v��^� ^��.n�����om�!�J:O�m|�V�kw녲�R���`G�{I8wг!j�fe�xqG��Y�Og�-���⯓s����>�P���:����T9�Ykhi�ËD�r
����g_������p�>Kä�@,���0��P���?��.�߮�E�󖡝)"VMQ�f�D���B�j�|7�}���>\DP�`�{�3��-C��]�ZU#x%���1���󼚈��4��2����HĤ�ݬ��4*���,�^#���m�����)ȀBk~	$���� qy�9-�r�&��]���x��t�sk#��C�츆�T]]�B�!�d�a�n�`%,��Q��'D� ���B��������<�/XMXY8��Y���%Y�򻷀ŭ�2#��eޜ�B�����@����_Нf)&{�+�A\Z��E�ѱV�����ʼ�g:B��`�U�wgW�K���T�3D]�	!�U���/�u �WI/6��7P�I��0���	�ʇ�&<�+��YO��N���#��:T��x���/1��֣�����~�,��IԈ�U	;:a��zi�-7	�=�<jR�>�F'"몥�s5�b�-�1���A�y� ��x�~J7�&G	�s�ɯ�lO�a|;Ԏqƀ	�`�r�g��Ѧ��n}�tNd�!�-)�;�`�����U�&KJ��8Q~�s�eL�Y�%!(BCF������B�{�ZG�z"���ya��I���}x�g��8�'t��+��h��\JO|��-����7>|l�-w��X��r� ����׺����q���AIvk�~�"�<�Ԫ��J:����QuXZCv�r���<Uw��I���@��v(&����/��(M��߄��FWW�pA��#�v�Q��{(����h[�_�L~�1�݌�jd������
���R�ϙ�T�h�΢��yNC*Y���M7�ɘ�T����h�iI7k��� ������Y=��e��2>^��&c����B�t8)�*�� Z6�8��!����r���3ߋ��Qv� ��_�jS�� !yuC���;�#����M�\�%� �^�S|��xP����{O<dl���ة���c嬪���eŷtE��M����e�H��ܷb2��y��Z�������G;�*"�4)Gq�!���4�d
	|Mr�B�b
�̑*
Q����kH�!�݁&�Z%&��k����Ct��H�&$�w��_u��#=�[���i=�hax���U��ua�x㐧\w����N��K�b�r��A��`T(��'!4L��c��D��D���J�7�g��`x���HErC�����qye$�o@��_�;W��[�_�~��^���u�؋�)j|��K�c�e����">�����b�:�LGbH뾶�$�nO�g-�˻`�E�0���n;w1S�`�C�{$%O!����uȽ{��� ��O�TV�Џ�U���Ex���xpI7�Z���De�u���
����
2�cj��R��u.uyy�R����e���
L�FJ�J�3ޡ[ �Z^u?A�u:�ڏn�i��Pb�S&^���\�P�a��؜F�EA[H3k�ɻ�%�3�c�Pʁ����j��9��W��-�D�kb8@�C��:|���b�vE�L�ۭ5�sY�Ė�ױf���/��3��-�t7�A��k�Ҍr.��0�^��L�F�.rq��uh�ۉ���3q�����̙Y�d��BPY�] �m?�ee=�"�(��:������/�<~L(d�P_�ģ��c�}�ӣv�(�ظ�EF�k��=�T�"Y��,��Y�T�h�Dn;���f���6���1��C��� �#�	Vh�>Y����.�q� �r�������`^իnr�4#�Z��h�!]|��'���X�"��2e�ܾ~��|�l�[�����
,d�T��:^�8uĝه��<m�|t�NH"?OD ��ZߚdRy�
��=��J������{.ۍiڴC֗nv~�{ƆFzadiq��^�pjui�$Ϫn~6E�ıq��FA�i�0���&x=3��i���=X��e4�w���p�.�J�[3�5�ϵ�=QBi5a��C*hօ�5"᜼���l'�F�0C���媌HPO�#4զ�Rϣ���X���쳏M�u,d���Qr���=�-�K��U9����٦�v�v;�3?D㙓�^J�5��Q�6���˸[և#{�R���٣�/FK�J^���cKp,���g���\K�yI�;�z�C`�0�xté(����ՑQ�� ���e\��e�WoSZ�
�����H��z���*���ac	���S�7Op�_���r��>�VPBA~L3=��w@�.�慵�x�~��?�q��z���� ;���'��ć\�c1Dφ@מ&�����N�=��|���u�2�������i����a�Q-���̯�]�F�ݛ�u�q�iX^wmaE�j�eF\��+SŮɦ��C��F������Qt�����*_��z^��1����;��e=FN�7i�Vj���wB�=8xzBx��� ����1���e��$�mi9�	