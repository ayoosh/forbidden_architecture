XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u�A:a�j��a�W;�֔p��{����-����?���Ĕ��vd �R[ �N.SK��ߣ�4�h`��Wb8��5Mb�r9q�]W�	"�j9g
�'��s�,sNl#��Qu/���o"\[䀦o$FalSγ�e �qʈ���Y��{Ym�?�ŵ�eo(���֕b�`Lk�Ne]P�\�����.���p�
;��+��Gv�	y�2������=�\�Ư"���\��v%K+���U��������	"5�}�q\���LI�v��oL��mJ�r {�{�]�������bs��&�ͯF�pK	����B�bX�����n,������E���&L	2B��3R��:1ViZ��鵦�I�nU�a��Wq4W=9�5w$�۫�޴vp�P�+��C� �1���,hl���+���GO�%�dL�͛`�����'4NU���������s#�ʑZ����G�m�?HG���ގѬ�f��E����T�rF��p~eظ��3��>�$.O���eX�ڱ�"mz�M�>�99x��x!�ֲVc�&c��?��R�_�*n��3��Pk;K�34)�Փ:�7�v�~"'�%/�󼖌>�Q���a�K�x�<�K|�>R�S����x���������ҥu}f�4���sQ���o(tB���c�r)f`�G%@^��?"�Œ��M�$K�SsB����*Zf��<��D ٻ]]�ʜ�*+|����Gsit�c�(O%x�#�K2^2�QQ,th���Oؐ����XlxVHYEB    fa00    2260��+YS5��q!�Y���G'���/�J�́�]���s����t���<�~�Y%��;ԯ�v��җ�����`�u������}�޵����vs�1�� ��J,A�~��7]�!�pm,� V�3��?7�ȋ�l�@�pZqyZ-X$a��+ ��,e��ݜ�VT�b.�~~K@��EˡБ/ ���qp��2�?A����b�9����U?�1��4�BȺ�����nrN�:��M{ʇ8/�@Y�����K��(r?(c<����`m_7v^���2f���h�\���}��^0�.��h� �#�r���9��t��X�6'F�f^��W/����X�'�w�O&�eLx i�hꘞe)Ih�[ƝNkC?�sTD!��a�h~��<X(`'C��]d;o����R�E��7Z�^:�>��qUn�Ee�?Gae?��80��<J+�)?���1�T=`>��S��$�ib����{.jP�ZvB�>O��]�W�u�̧4-!�� ���7�8���K�#��?�/i�K��w�ub4��K�X�*�Bյ���Z�2��1�ۣR`������<3B��F=���J@�+H��c�4=@'��Z����*�Qvo[�H��}&	o}�BM��2�.j�pH����oA�����еkb�0Rj��$|�/c���LUD~ી.%��Qf�����\N��z���mq�:������㽆_+zj)�S����}��`$ܔ7q���Ǩ?��%%��٣�wsعi����<��J�=��k��O�JRd��}����'�~B����ɒ����j�	�b燲�$�e��c�烊wMZ� ��N4O7����e�}����,V�g&��k.q2-�͐�Ց�vӱd5�����8qsf
�Y�k�>o�Я6��FԔ��BS���1H���k ҷ�L�pXpE�͔u���I��\��j�єu��1�=��-D2��uO�"���0�<:(!�(}qz������c<��BQ�ZŚ��W1���}�`�k��׎d�j��@��$�uZ`��z��G�T�};�ƪ��?	�w��$��T��� �	���2M�f�_�%��F��:�r�v�e42�v�Zv�N�X#hU��>�L�R��֗��üU�=j����V�~|xpO� SDK>��Ih柴g}K�;��:9oI'� 	y�
�{��K�C�<ޘ'4�6#�|f����,�t��ͬB�oWB��;�m/o��sJ��ݣ��H��W�.)}��C�Ϳ{�a����÷��>�Kn��]��e:�����j��Q4��U���	^��v�f�U�C���vK�����y	�0ŕ<����A{p�	v�F�:�*���ې�t�(�10t�
~�i��X���7Y��l�{Hz��W�p��-�J�z����k��ޑ5����@16�yw�s���˰�,���I>|*ܢV��n;VJy5_����((�g秙9�Z4��:q�(4�tf����-�P ��kN�Zs�,K�W/��z��Ωe��˛��O��� ]4[}p=�B���^9�u�Y��iL�L��H	҇����4���	+���8q��f��Ր��O�۲-	`ߧh���<@Udn��I�'��|��>x���4�a,����{�P��e�7��R�*�0�}����O�W|���B�BS	o)�H#.d`F�ﰮ_�m"���,���zyÛzPذqY4܍���V�����Mk�W�׋�ރx��M��E-���OČ�*$	e�{S9���8SU��H,p �ՖC�ϫ�NV����G���� 5|�#���l*i�'��(�G'HZ o�	У�5l�+fsb���a22���/�/,�8�3'��7�H1���k\R�d�~a)6��YO��m?��O-��׹����������G_d�e��q�)��e�����0�xZ�`������ܶ�)ԄH��x]9�kE�
C�5X�{�_?D�%���O]�Y@�t���f���~���ـ����s�]�>�?2N@�NG���N8�T��%���Q�s�xu'���{�%9R������ZQ�M݅;Wm���hA&!�
����,�g7�몬������D�Vq�*�YHc�-◰g>�/jo`��L�ihB!��/�j	>�M=K�Wy$.Z���bi甪ᲇ`�@��=#G1L!�B�w��<a�"����p��x6��ۡb���D�<�b���(�Z���]���SLR���T|+���>������x���8w����jY�V�f�g�>�3Ǟd�URs���]׮�6���5�H6LNRѳ����a�h&H		*T��L�qnxA�KX�/�/&ё��/�QǏ��ؒ��LW7�*v���n���m�b9����TJ�n��<w�l�=G�<>�	��fȰ�����Ϸ���n#P���>͎����rxH��֖���Vo��  ��l���N)w��%��h�!"�l)b� ��8�w�J��ˢ��8$�6�w=H|N���%� ~۹B�,N��"���𲃪��Y����oҬ�
ȳe�k[#So��X�О�$&'������7;���g���cU�4���=���،�Q��t2+� 3;����|{$B�$8IA���֠�������5�tZI�?�G:<����G���r/wҌT�
פ%�.�Ц���߷GLy_	�@��87���c@R&��m �ל��� ��b*HN�/�"�\�?hO����`L`�SW��$.,S�rʄM�#Eq5J��G��5V4N�7���/�G�9T�K�Ο���H4$퇫��=�3l�P��ߑ�%0fg�)ռ�e�[[@B������_<�.B�I����ϯ��i\��h!����;�HK�_i���R]��L��&D�E���%���a��_mR׫�pp��s,�} r����bJ�!a���S�"�Q��z��L��ѡDS�$2��S�q
c�$z`Q��)�!�/2>�!BG3��~Φf�uI��(��f��nE~��S�޹�w��7<��JO�{�y"��Q�[u3@����Yxo�2~s��D�S!���V͑�8�r�qt�78�C�	�0�!��Rc�[	�dYz�$3���6q�	9���|#��k��5p
<�hn]���+/3h�����v?�g��mh�N�s�ɀ���;"p�pO��E1n�����;S��ξ��-���#=TS����k��:C��*��W9�ESJ�����Q��۾T6�v+|���ɶ��@�}���k�dfͱ�����dZ�0F_����W�y$L ���=ʏ���R�:��n�	d��YS�{�Bͤ~�N�����3I=���h��f�$�I��l��8�\��9/�� g�|Y��s@��^6�}jF���5��h]��7��뚩�U|��q-�M��j�Q�ʭ�L���g)9��Y�n'��$�8�.�!�J����
/H-K�]������͢�L��(>p�յw0����	��8"&�2��"B����^:���w�����)��*v(}g&�,[��^$*c��ݧӴ?|bO��2V����ؐ�be22�ʰړ��&]���G���'rv��O��~8Yw���=�&D�xni�D)L*�H���(�Ḟ��F�hi��^ϋ�O�f��z���lOf�@�G��@D2�v��vE3��d�� K�޲K�[�'����2%��Q_F~$����(�5!��㛥����n��$���K��]�泃u5!`�.���>/!y����;��LF͐��Y�)���Cʮ��X&���96
�r�n� [�/-��W��Y��is��Prh�c"�NT���'^�z�#	_R#S-�����FDk���մ5��/Ԛ���^u%JoJ�a~*��Y9���>ϩ���`�p`���S�$~�㞨�Oy��%T���d��S�Tq�:�7=�Poe}�C��6(���ޟuL8|A{%�J惷Ed��z#/Ҫ��{�fl��(�S�Cٴ�I�<�QOa�q�:�|+�v�k9A����GL�?M�B�P6m&?�G��Qؙc@1�tDAyn�����S�"6QgXv�%>�#ߧ������ X�U���%޳�H�v_q�ᐛ�jĳk���?M�x�&�<w:�y��ڦ����s�|�*shA���n�[#Z"��=��H}-���kML��CV�>X���ƚ�U�I�<%��>�<�d����<�鋆�l�fs��u*�)Φ����Z`
�p���s?��Ԯ�%n��1����a�8�k��'�R��O��lų2?f�	��C	��ǕNfT3X�P@P�|�y��g���X����8O`�;����|�4@|�uǛq�3�c9���թ�J��!���ɡ�Y:�\���h��Ů�O��� 4��Z�1�qDO�q���X�ta�v���3~�*i���+���H��\�$��f.�������[q���&DK�@���m>�N��Er�U?6>ہ��Кl��7"F>������Lx>F���^�%V�mP��7̛Pƶ^�[e�k��PɊzL	�:��9^+-�:�T���s���O����2�w�`�*��S^�~�Fhs���T&���-�)���ο�>�B��?��Q�EgPO�>����L��s��Q�Åt�P��5|
Q�Cc��{��y��(e>����#^\ꢦ�����`���٦���;!@���-��S�Jj`;0�o�z�Œ$kG���qq2�A��8y/�K&a��9͎��˞�O�h
آiW���iΐ?oq#�������6�&Íu�� ����|� ���;�"y��8@� �{���ǭ�іC��âX�e�bsO˂�E����'����.$w���"�1� K^���յ�
!�v��~�%Zw�֧=�i�Ɯ���rg#�f|��$�g�S�a�[T΍m2�@��c�=�a�	�� c��
�x���턺�~@_!�X	�~!&-L��aߵ;7�S`?�(vx���߹�.I�u[��-,`з\�-��Q�f1Gw�q�_#E)zqW �g���I$�,U]&5z�F!�nx���+ �@�#Bg#���J'��E#�,b���Wo�d�V�U�Ջ���6��D���Z":�����������b]��pY�H�>e�������}�)&�Bd[���>�B�7z���M+�a�L<'J��c��X�TW�|]�	�Ń\$y��ҵ��Nxp��I6
����BP%������������%h&ɐs(\�2Z���)A|��A%��\���Ū���J�&{3�6J��U庂̫@ �[xc1*,�������6
ݜ ��KW
��AZ1��IA�R���{k�d��e�Z����U.�<��b�V�6MjD�g�VL����}�HaJ�i���n�:�Ѻ}�^_�Bը�MiWm�>%��K'2P�Z���%ѝ���T
g�&u���2P~ Ҳ9�r�Ո�$�(�b�t�%������uS�|ˮ�.�e�qL]����S$��A:������c�8�1X�5����=���� �*gK/F
[?�R0��U�6��Z��}��h�Y8'E�l	]ؠ�c�|K�+γV\Y�r5��4����b���/�?�M���$�I'��䇛'Ld�5R�p �g����Pߩ&
�����$G�-ζU��MB�?r��'X�+׌9/L��B��R5�QQ���,��]�T|���jy$�&sU+%���%����OAMI��\5�mh#��
�U�|N���`�v��y��Ћ��脨t�dIK��&	�Qۙ����2m�cs��r�т^��Hs�.1�_iފ��q��x܄��]j��~�� ����n��@����8~��X������\�+��f&	�J��m��λ�v���L_��/v�����v�����4uF3�0�$5�K�[��&���G!�~環'�c��#kwQw#��B�P��\�ш,�uxy��/=>@+�j�#i"��ߙM���35�+�*���9'�:t�QZyd�AR۽$��LO@��w��%��*�{3��o���6K��zh�W�[�E�j��u�N�4hG�h�@!�w�w�.��	�**����d����_uC���G�˭R�'"�`Y�;���p�{.C��M��UO��m��%khV��r�jS��p�L�[S8X�)gRb*q�7��"�E� ز�T�����R��7�������v���@j@�o�W����ݣ��=�!;4�NK�j����~NA6����]��^i'�$�0��)]��N����O�Q��9�D^scI;��v=�L\��a��0�c׭����lMM�ے��e}���b�U�����;E��Hx@�Ͳ���=Y�1m��'���J�ʎ -%��������� �MT�Q�2��u���B��r]D�A�n��um"�g�?H��%zkt��h:#ϡ�������vk<� ��1XEM�A@�iR<��~�̧n�t�U�֛��y�o�E��}���B�Q�j*؞�g"ᲁ�tz�� ��5�Lp��}`�K�e���S�qʎ�
z�,�����Ռ.1�8�5WQm�º�����^�^9hL?�Y7�"��@�J��VV8 "���k c'���� �!teM�uG�k��A
7�����W��m�M���:���lLt�BQS\� ;��T�������!��啯>lV�Y���ʧ[����s<��Ӆ���ƕワP�%|�}�Z��{��\ں�j����`�B	Q�v|���ZKe���1ӼD���̩�]-�i#��%v���Mٟ�.˳�>�A�������p��囐i��K���<�phi�+\�5��9�E��{%�V�P!X�E>D�T���$�Z���3sX�DRЪPn({��!c�iD�l9o�����2'�/ƄZ
�=��ݫ����l�f�ߕ�%6���B�@�<-�d�o
ŁkX����B�yvA[9ƙ��$���Δ�`aH��l��q�4�t"+1�b��&Ӹͷd��j���횈+��14(�4,=Z�[ɸxupVt��S��/�k��OD1�t��#���#���4q�����"���9�H�D��-�v!>j���mÎ���G�io����1'Pk��7@���
�ڒ���ᒾFu�{��'�����%3L���GB
ڣɉ�9��&�u��V��d�!�S `�MU��<�UA`	3\�<vj�`����\Y�V`�7tn'�7/�s12ڢ_�6#CB4��7e)ӑ�ͻ��
�m��n2���yUkc^��u�x�<tO+��K��*7�
�zs�(^s�9e���}��5�"�b����C����K�����˲_�:�og�"���2X�^��g�c�G$X��[��b\<y�����@i17�+ަ�ήϋK$�+�������9�v�(����hw)��i��p�h��K�	��mC7����=
�8:y~V�"?��#�@�y?��h ��hes�_p�����0��2o�b��%ٔ�<�9Q��#����i�3���?9�c�i"�� �)?�"!�w����s0;;K��0�����$Ґ��ɐ7����)ʼ,��Y4^=�'_���t�x���Jf1�����]�g��r.�l�����>�M0���̈'c��t�r�_9��C�y��6)b�
L�G�#~H��6`���T��6$����l��M�06�T��?�v���Mc��'�}6`��)�r	iFD[6��OhN�+:>�����b[�<�U��H�) �>n�C��b}�r��Z>c8��d�I�+ǭtf_��k�I�5���	�Q q~���(૽�(�4�����R�	&Bx'���pk��&-v��7����	2룐�Ʃ�wl���gcވ�.�=�u 6hj��ʵGl��%r-��"�O��A��8g�g����N�e�5�E}��[��V|��E����Ru`r���"��B#�K>	?��r ɡ�!
[<�I$��+_{��r�(��L����#w�^{���N^��E(?��݂�}�"�� ��!��l�"��	=[>7Kwտg���<���l���ud�&i"�pw|�gVn����s:�F{@s"��U�$��/���O3J�60�}��F%�5�/O"��a�ʄ6q���9 ��.���o =��c{�+a�����oX��=�0a<��v+�l^�r�	1k�a��س.mh�̕%���]�2���Fβ��-뀡D�#�����y(�n �a6E���ߔid@��f��;,��_�f���n^��[fKR�<���?��2HC��p���;���Z��x_!�h���=��������{^vK3 �f�V!�n�w}_�`�s��D�$8��-��٩-�,DK���)�Ր�Y�ߞ��u(�D�;��K�|Z�A��r��m���9
��`��&���%h߁o�Lc9Y�q��F��]�4V�"��)8|�|R���\� xA^5Ĭ��x���m�}��[YG�8���s���D�3��: t��w4���	��U�j8�\:�g��wB�[�m�Pi|�ث"�22a�0I`h�D�!�5����sR^��K8��-�'#�w!�c��.�\3*����4���/��-�&E��)݉f+Xnt�Ï�Uu_������ŵb3Q��f�']T�*P���h5L$��v��m�SV{a7SXlxVHYEB    674c     5c0���1���E��>9�����{	�xc!�,�U���	I}h!IxfF�}P�h݆H�:L��8��J���;�y�X�}Ҍ=$��'B!�i����&1����y��cxL���������[�����E�NT�
9j��9Vx�f�?7�����pP�`i��L+�(9��W����v��S�.��q�]����D������>�������yʚ:I-7;���(����ݮ��߳"h<I�n�K�0�����2��Ť�`"2}������/���hg�צp�Res�=O��IjJ�$!m݈r�tX}I��C�pL�+�:;�Jl7LL��8�.��?�Ĩܛ$LVo�J�G2^�\���_��_��dF���?�sI:���n=�x�s'�:���Ôc��h��)h�x/w]��$D��>�DÙ�>��Б�u�tys3�,��#���~�I�m�x��]ZkE�!B�r�Y��	"�\KEsU�t	��^FifZ%N����$�<BW��X��h%܏R�:r��=g����
}$��=,vR�����v�0� ��V Q����0��L���}F1��X)��4�z�H�Խ��L���&5V�/P,�,���y�ѕ:[�~�`f|S`CU�V���[(4��G�պ��������"`?#\�v�co,.<~"�W~���]� ��?^WΙɑ��󑟥��˒S!��*E[������S��@JJܵ����&�A�ko�?|s*�ٞ||�£���
�2�WĘ��"���^�T��'��8��S����
Q�-6���e�Q���+����W���>ٮ6�i�_���E�'#��j��fp!"?|�"x��v��+xwM8oK�6�_Y�C�d�j�iL�Q���Y��mPdW]�Æ�ŬAn��0�f�ԃ�&ML��Ғ����U��wՅNB|�qNY �o 2JH:��V�nDA'�KV2��"H�ka�]��P=�?o77��H����`_��𿐎��R:ߊ�E&p�����c�z	r�,�=�_P�ÍJW�;<�Z6"�-�{��i웰�8{)���������彈���&�_��
����(��Gi�k-{�Ϯ?5L�a����h������ʗ������֢Z�g���CJ�����-�~BO�!d@,LX��D��������G���`o9s:Ǭ���g0-��mk��,0WְϽ�C��f��@+F�a˥J��"�5�:����Ba�P9E?�ڿ�^ӱ$XS-=�'U'��;�PH7]d'}�ߖ�L?����,M�;<D�u�:%vg�����;]�
yL��R�bJy��k�(���/�a��Ԙ�$ߌg����ΑB�� �[]��_Io/�f�ļ��k�V� �sU���krᩤ�j��kp�u}pR0�G�/J�d���t��Ֆx#��O�W[A����[�� �@&E@Of