XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2�DǟR�CI�w0�&//�s�'{��aҙ5
�W[����NQ]=�׀,�u�vy�vf�:���'F�x`�m�OX���
u�f�4���\�:�;� D�`�H�"�R#�@�hZ�3$%�����1���6H�GE:�ws�\2?v���EЉK��0P�}��>�fv����
�I���"bg��m��rĶ�[4n�ިB,������� �՜�M��¼�b~3�fCT���(H�i��]����,����hZ��F1tec.��Ur��-j˳,*��A;�Q�����c�'�ЕS�w�G��Q3V���=�"0r�j����I/L]_����y=^�.MB�.�s�Lh-�N>��$T᳦���KKƪ,d_x��}}�#B�WLZN�31������W�;�����h�xH��	<o�S����oE�-�`��[D ��u����"�7^��DP�jV�x��JF&�-]�/UޞoԀ� /'��YaAӚU��"B����Ey��4T/ 5.o��t�c%�r�l�O{���Ќ��kk�����p�؛e��Qj�>}�E�y#��M>�"`<�l����p߇�zH�;q���c����.�����������=��޿q��^6.��-��m�C|�?O^�#�x�P�����dv���嚲N�����jS<'�J�4H��7�%��4�^붿�o'=ńK2���i���2�`#������)�#>���h�O����.���VN7Η����~�l�?V��?� ���c��g]XlxVHYEB    5cba    10c0kJ�b�;�d�S�T�\a��k[��*��c��i�ŉ4���(�rS#����orx䉝�?�[�*���5��ˏ쑉)41�C�t@�ˊ�yD� ���[Xf��L�}aɋ�<�}�c/�:����n�J�~�nV@&x��c�5�����y�Ӣڲ<��.Z�4ّF�0#j<��Ӛ<r��'���5Q�e�Eed��Gc���;�Љ������7谪�YU�o��2�k�o�Y��>�'$�O�\��.T���q(z\Ο��[bJO�x
`�T�CV4�m��6�TQ�$�#����tV�92-���oj؟1�����h���}C]�����-�+�����\*H�@v��ņ`�����K�i۝ɨ�[ۨf��4�G*�]n�Cg�a����5i��b!�e�o�\=Np4��s�S��$Ȅ$v��F�ձ�l$)	w\.NR�~�
��s�b�[H'���12��uZ���߅�Ҍ�inDK@N�R�<��u�Q-��2�}�Ly��['{��LF(������v�b��п��ru�b1��a����:�t�O��t��G� ���wtK�[��h���5��0 �uQ�)+�_(����hǃ��͔�3���wO�  B��8�{@�،�32������P���A�3I�ц��Tc��c�V���fߋ"�\A� %x/hه�7��<��g1�/��q�ϧ<:���&ac�R(�;�O ����yG���޼�!Rz|ϋQ`f�<;8�U/Q% �;m"g�[���b{�+����|1���'�I��L��� �P]���&�a�G!�G/�J���o߆�zFפ�++�_B.V'5�^�납�z\U�Y+�m�9�9�vo�B��x:�6Q�+V��KF%�77��	�hS�Oqiz���@�?F�"�*aR�v��R��k
Ě���Ƌ �K렩���y�X��-�58PD���Ta�E�=s�`������K!�q�!s���%�
O#.�S9M2��su��*��͑�d��O�m)r{*o��%�OdA�|X���&���җz��E��ۃ4V�)z��ex	�i@������J>>�v=Q�s>�棅��Z�Y�h�敹#*^��;r|�dw���e�_ �f4�a��h��Գ)����4SE�s7)��:� �f5��O�QU/	xko�̖g��ˎ|�φ�r�Cӯj`�_����'�>B�u��ٶ�R�#r�=��Y7zO3�Jov���d�%�_�cx�a~��D0hɘ�	�כޛ�X���|�����Ԑ�8
I?���z����-ª�h�R��v��Ư09�|��M$�i��?�F����O���������<DS��Y^��/N�ֵ���w�-���i�����Q�u�5̮͆��FpH�z�;��Ĝ#��B��Xpm�2DW�]̥1�	��G��g��9�����C4���3��Z wz�I�x���̦m�lF;hǰL;����0����c���d�BX�@%	�j��)5��V��!���tt���3�?A�rI�s��P�ɶ��[���z#�6���r�sS��������U8��o��ƿ���<81>�M)�n�+!x�ftڀM.8��#���G>��������}��!n���+�cڲe�tT<�]R�l�r�V�=Q�CQ�3�~-$^t�G�V��子r�B���~lK+<�gw���E>��}x��j���T0+�7�(�m�0����I�7��U�Nh��>�W�#�|7d��Y1�(���+!D=�'b4��<�y��p�ѓ��q緃�r�\<P=w��>k�q����w��tŪB6�,%���;�S�3��*W�P�\R7VR���K:���:��P̩ (uY.'�O�s�|8Ck?�^Z���y�yY[����`�w�#�o�!�"�H�4-����'Bj @��I�:�z.�[��hB��2x(4� wdzw������v�,�����T����o��<�y1�n�8/šg��3hmK,�m�((���`�_�)[���'bLR��\�=�/��?Wo1���}^���{@�@e�O�Ӱ�[�.=v�0�*���c)�EЇ�2��_��DR��# 4����������X��H���y_vB3�^oB��x=?��tJ�R{��0L��i$#����2E�o���h �C�1"3�L�ߢ�"����軡$)��h`cs8�3@��~I[Y��m���ߴ�Z��9,��)3��F�*\ߺT�̟����(UA��۸_����Fz�x/�P!��f��-5qt=:U.���f��t�Px@�uC
�-�sɦ�OP�@ٳX�Y�Y{� ��k�5�����
�-���Q����{�΍ ����)�2S	P5���"o���X�{�F#����CX��(�đ+�����ʺ��;L��]�h[����?��	>�� w���{էQ�r,+
��z��BB�'�1�}WY8��+S�-|���U)��̡�7��//IcA��/eEf��Y�f��:�1�i��$&]��8ym�u�$P���ǲ���dG,�c][rX뾫����;���'׷2x?�@��ө�Z�Lȳ�hSBE;��c��&ߢ&�:~>)�K�v�m-״�o2]	�wvD!�26!��,X�[���A�!���ma�|���� ������ϗ������4F���x��;K�oȬ&qN�)�6��e�x� �qp�;5� �PiZc�Ž9�R�:n�6y��z
����o��dw�OW�ቸ5��yR�$Ht�_�KԆE�%��?���-�]�i��>���,�E�础����ȋ+w�:�g�(]<y:
l�̎��ÊX��*�&�����(.��EI��'�k�X��+�ю��%���������E��Z0#��K��R��ٰ}xZ�H j%Ycxvͻ�s)���x��P�NE�����r�t �HZ����iwo����ڬڂ�m�d#ـ=ƈ��NП^�`��D����;Pl��Iok|�\
;��緮�1L���󬯨8���<m�wKR.�x��|kH�IR$�4�D'C�B(���<pA�l
V���{�d�ן�|K��hv�	�qi�����Bz���U �V��$�AϏ6��6Av�|�U����&%2KS��u�y�7 �u"*���Bo	��v�$�M�A��L�upq�&ǎ�7�p��Q�	�Qx�-} ���Y������d�g����[���VՍT1���o����S2#�b*G�9㱽�x�������7��GHX��wG��;p�s�+��!0K��j(�_���\�;E]䱃:�ʮ��IQ˭��ck�\y���A[�M��;R�ȂUs�d��*�n�}C�0 㵄7�$��
)l�!���Pa��q��l�9���J���1l�*ķ;���4���c.����=���Y�ף�����s׸d������ߜ��o��O�7�0
L�B���p&�W��˼�MX��g;^g{�Ӹ��f�֌�j��Ǻ�g��)~`��++w�䓁�qcĘ��}�mR���	�����ru��i��dO����G�� �t1k���C~,�q��BYEʻI&D�)RJ��,}��ăJ�Ʌq���Y��Ro%O�R�j����۠y��|r���m�`g�q�b��%��oh�˧�[!n�pg3�LV��A�9] ?Q�0ã�)�ƪޖjɋd��t^"m"���S�a޹"���&ꃨB�*� r��^�Y����Q�%�hM�y* ���[��^��l-oG���c�� ���&V���#� ��h���[.���3­C�������B�;:�*�l�8���;O�*��:�2_���!�[�?�
��:>�TS hn�!0��|���#@f�d��6l��)���!sh��{$���y��^�[	хvk���:%ڄ ��2=[1�|��V�xM~��)}��D|�W-��X�䬇;n�N�!#��J�ާ�5�("�fe��үA���a$~�H�'?��ZH�c.:�M�@�%�� u�
��Bd�GcP��A&��Ȭ����;<�]^�O&��4�ѡ��Y��8d@ܖ/��*+�����u�<�\$�)_��:��/o���9$�u����v��x�$�B�x\r�$~jJh�
���D�cI��'��-"�*�V�S�t�"Q�D�>��w�,ie^ӿ$c޸@����>
����+�S]�I��/"'$ |5jo����8W9�H��:fml}@�-