XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v ���g�G7��Mk=HfP\ {�u��T�����ˣ���n���W�z!��s7t����H@�B�UCg����F�u����(�YHz�!3P	��-����q�4_��ˇa ��o2dQ�>��'�+V���d�]�x��Ba�v"j_�K���ZU�1�4���~�N�-��={D��!�s�T]t5��	Ne��';EO���5�Uq��YW��lT�=���w����О �@?N�x��f�s�g�,�+nF���S���v��6��uϗqpU�ɲM��	+��>[�/2�m!��#)h��m��BCEU��/����|����Ɔ(�o)J��b]��k 	i�Y�� $���eM�2�|���g��@��9�C��|y�X�VwӀ��S�`U^��Y�U�Δ۬��F�h�ԅ�p�%䕐�����qB�fx7Q��	_���ѧk�E=)d%a�d�[n�rI���\���Z�J��"�"y!j����H�+�(	-^$�Fj��8cy$얉�?�Z�����4��<�(��~BD���f��T˾���+/��b	�%�:�����b"����d��-�KT�B���\������qѓ�,R�cfّ��]�Y�G-Ŷ��
��[�W@pP� ��U��C,[�u��N9;�|��2,(ZΥ���vU\�R�r�p'�/BP�}h���e�|��r� Z�:���y����tH[�t���\���i��\_Q�8&~ƵS���K�G��B�l9��O�~�aʢXlxVHYEB    fa00    2020���5s޾|a�^�9x�.d�{�A<�O�\'̵���s�Y�N��T Q-؛;XT��˸��3���<�I�Φ;��e$��hcmb=��k:���kMi��}��]�;.��|�6�4X95_���=M��7ڳ�n-[�����pD*�L�M��?������`�uɇ1;��{�#:�*�>l���;M�ۂ��}E��VS�WO�0��AK,�ٛ�#S׉�)�@r��*�� ��5CN��et��O��v2�a�&c]63�*ƈnr��~�Q0��
���v?�����X��5@Ś��A/]PN)��Yھ/�b�!���c��jJ�0�MW��8�	/b��_!X�o�e>3L��?1��c�С5��h�eHS��L�ȷ[�� ֞��y�p�X�49O�5�A����B�.���-BB�����}��oR#9�EQ���4+�`Ϳ��^�'��h�{�*��Z�Ml����L����~��k6�l:L��	�=4	Z�.4C^삔�<�l����tl�A�Ι�Z���l�; /ĕ�0��徜 �`��Wx���%�1�����ig᝼a�G�Ϙ�t����x����ovY�MI+�=YFD�d�A}������R�7�n=�@&	���8����ѩM�
!��m��N�9��~kJ=�v���d� ���n�������;n����F#�u�y����)�y9��m��H$��!��U*�j��G��&�g�� (]��iX�_��(p���,�s������|���LpPJ�nI"�N3=u
cG=O��π��k~@R󇊲Z�$�@������m�h��qko? ��sGЧS_5��Ϯ�J���������Ǣ��%Tx����aw6E:@�ۜ��E٦i�y*&6�>�];����'g\�:/���ͦR/���o�j#�:8a�Ơ^[Zy��~���=�t��@�oDr�a��C/'�#3��`k��nx\Z܎R�9��� ^�E{<O
x���� ��dǾ7{��ߜ����_��i����뮶n�qE7��޳b֣���*k�9B��@6�F�g�
�t�X�GF�N�����>&���W�?�GM�x'IH[uFB�����&�6�uE��*!L�H�TͭOEQ���v���>�-�6����������:���q����������L��X�+U-���e�g���[W~k���*k�m.����ʇ���uy�'������Oj����'�d�P<�%����$�?�ݮ�D�Z�r����U�^A/�^6}$�G�bL(b�n�h��ֈ��,A�.w5z�ǚ�����Н���Ouz�B��aA����Yt�Ckv�1��d�P��d~*@Ș��^�{�Q�7o��냪D��̬ɨ)���>ۊ�|o׍�`���m�X:\j�a^F���]JM;	/�?b�R$�����̯�ں��{�Q�ӌ1�'����iڃ�л�[�ii��b�kI��%�މ�+�e��Q��35�@re�Cz���M�4��k+�S��������Bu�a⠇ݳ}�ʄNI�Kg)�k!���Qu���1s�{U�t�U�<���9,���mxF���}�x�)W�S)'��ܧ]�oa�Rbzx���ʳ��΂(���D8�7�/�VJ�Տ�����bt��p|�B
�6��h"
��r���4���E.����W��a{7��Zx�,�2���<�{��ɍ��E8����$t��[��Qg�_�9i4��欹�)^i�[x�	%%�uC�uY��=��2}�hj����������[E,�2gS�"������."�˛�L4�5[�a�f�1�V��=�);y�Q���*k����q8�7  ���IYB��~�z���1(�y��uߢ�G���fҘ{�ܟ�t����RgY�\�ԡ0���M�g��ޟ��'�qSGw0�7W
J����C:l릺��{bwgN�C!%h_�:JU�17iN�u�-G�z��1�f:� dM����k�̤���0��b�������b�&����:#�=0b�`O�G�gZ1vl�.��Rmɰ��� ə^eF��]P#�q�/�A�t_�dq��l&��98|�<��|^(�n���53V�^���z�b"2���7�=t�I�E�u&�X�L-	��kw/i���BTJ��Tm�������^	��K�`2G9��>�Ċ��N�X�V�z
�A����;��F���\�"xԑ���'�J4�Zp��d��/�ԡ!�^2���ez�nIX�+�#��L��aue��C��&F����7I��yM:�w=?��ϡ�S�R�_�������~U57���f����E���e��w�͏��O:����i���4�/�m��`�<�-4����WB��-a$�G=6�H	�[���C�HR/�p������W1��{J�ɐ�����'������o홺j��P�]���8�v/> z@���* ®�?<�lR� ����4}�M��B/��7ۺ�,i�&jדƊI.��Lz�#irN���Gh�x6�a��#�����6���!�S����p�|n������PV���!2��N� �Ү�@P��\P���p�N��*%�1�$6���5T�4EHu�Oi���������d����<egH�c�v��&������=fSq�.Sn�9oU�Wt��@�.�)@|�������y6�7�ɟ�t�Sg+[�R7��\�� /�������\R'�/�᝚n� ��57�3.g�Z{�}:�8����6JYe&+�A�:5��.奈]��^��7�����1��S��ҟO�[g��"�9o�K �A`��j]}��7*�Gs:�i^���	q�q5)pd��}����g$��A�s5�����8�4/ݠR�"L4uq��6n��Heށ(�"0�lI~{�[� ������~�ٚ^@�=��ymd�\���ԲO#x�v��<�q(�gΧ�C$����$�E�"u�lv�~��/� �(^o���2�Ml��;���Ec�RG8m4�qv�g���p�2k�����9��Ђ# �� �$��1@�Rk��S*~Ɉi�Pޯ����C��O�J�u=��N��M��r�:)�;(ݙb?�SsQ��DA��tR����.4N���p��{Tk���gO�g�]=�3ɚ�x E���}���bf���t�2n�~Q���^����[����m�`峕 �w��vq����C� ���&����L҃W�si���������kpG�*:�R-��Q�.��L)�G��<������Di��+W� �>��&͟X$����d��s{x������������D@=\kw���K~�`�C'cQ����}��P��7͝�F���}� t��{��U��j���.�1O��V6S�Ҽӡ\�Y��|�V>���6v�k��Z��/2ʓ�5m�zS꯬vT�2�v�Zc;[[���J�V�xuPp`-#8�c��<c�;A�mT?�{��1KyV��h?+g@&U
��T�u��I����a�\�D���:��jzM�Lg2i?��}�&t�Uš�4C sN?�DxJ���r����/���ޓQT��R�~a�ؽ������p`��fT��g*�O��7l��x�0�.'h�&vSk�Lo�|Rԑ���^=�IR�?~��+{�@=��5�`s~�vc/g��0,�xu���@�g`0�:���}&�pF!J��?�lf�k��|b�r��5`pL{������.`�T��c��gD����K��>B��r���Z�?:�d�5�_�_�>�9��0�Z��AXgNpz̲��x���:��r�|�J1�^V-z��:tu6�G�-JEe _���w�T�L���r""d?K�پQ��E]��8�'�}9g5��s�m�Hs��+���g����%�H�Aï�9�b��)��wF!���1[5�$�'tnKv�v�
@�6>��LΡj��v+~�r����$�w^+�����R�s��ϼ�n`sh�}}��ws!VKعh�j�~`+�iw� c9�ȸ����L�V�Μ���V�0�}�`Z�n?��g@�Ծ�N]��[�T�Lh�Ϭ��[|v�a�iM%��B����"� �����&���8;ʛ��6�-�A�vp����r#�T3TI��K�Ø�����[�W�	\�/��T?#�OC�7Z�����c�<
֠��?�d�Dƪ�_:�۵���G����nZ��G��ˉuԂ2���TQ�STl<�5��*C�[���H&��k�v ]�0�8�R�g���-L�49G
�jN���P�^�7�*���ge�� ����RR��Lb*-BDn�ѳ�ъy�hЅ��`� V�	TN�o�&�mt�&β�߷�-�9f1])
��E���}��<�\�a���3�8K��)*�m�x��]IV;7��Q_�$�jOζHٶ�j,6
�����2��ݥErS%b�sy���Kڂ9qp�y	�9�&�6t�g�9�;0Q�`ٱ�ֈ��
 �u�'�Z��V����j�=phtrm�bk[���5@6�/G��=�i�*p@q����Ťpx��;�� ��� ?�@�a���ó� 0�{f�.�k���E���ja���O�(F6 ,2�Z�1iAn`M`U���uQ��<}��7�'D��Z��X��K>�S����N2�Ҳ	���ʜ��.���?�r��ቭ��6��Ȣ���ΆlY�AdbliU�e��Q?�U���K�g"���-8o&�Z��e-�>Gv���0�_&��k6u���d�2����^T%#�y����@O��-H@ si2���d3G�S/܃�ռ���1����`��g�d�QXL��V��XEI�>:f �z�C�o�%j��r+���K�j�!�)�Ά���,�Z
H� �O����
ϧw�4�X��$T��"j��^�~�J�o���a�"��,e������y��t�uͧC*'��`B��[k�#��f�οd� pB8������*x��/��~I�"��=����� ���X>�Ѽ�NU���=Z�lT�ٲ�y��N���/ڿ�CO�k�2��?��a�Bv\֖�`������7X1�[��!d�I����C�EБc�U8�Υ���t����8����B�����p-E~ī�f��B�X��(��b��� Tz@�pC����4��p��]���e��|	���\��K5z�?���"�"fa3��OY�su�\\�.Ke	풊���!{���żo*��&ԫ��CW|��Ɓ��3�u^=����j����Vx��RB��E��iqg�^&�`B\��"^����h-^����6���Ÿ�d'ň��Ec�FAj���#闀a�y�l�?�2��µ��LW�	���|ʙX�JY�,y��N��b��{�rNB��_OBA�0X�m[�	A�&�v�Ό06�����wЅ�#�Џ�����}Ǫ��n=m���Z�����~��Qcl%T�n2��󞄓f6�|y�6��x��~���p.���(n(V�o*���wWF;n^w�$N�\#�kA��1�"ǰZ��]�9��q�Cj�B?�M~�d�q��]�~����o� �<����LfX�g���)FUs��>㈑�{VӨ����0��Ry>'{Mm��ۅ詤����҄��������V��xn�#���0��)�s�@�:ZJv�Q�vH$}	�I}KC�2�_�_* ���d�P ��9c�P�V�ٽ]��Pk����I�D�B9|��~h�����7&Q��D�اo��i���Rj��Bj�US+ �?cs�F�:��;�Xb�8�R^��TT)����� _?Yɏ��+���g�H�x�|/DEe�(��o;��F���|=��o�x�Ӣ^�W����áϜ���I��%5k��t���J j��*�㇟����]��'�Z�,��,x �������0�l�av���#3D�5��2զ�� �7u�����9�R�~ =�&���w�3��&?���m�|��I��CO��I�v��0-�&Z�����w�<�$-f��U
jv�k��
���5OE��q�a](���6	��_IJ���2�j�-���$�&�U�:�Dz�������ޑt�4�ܚ1~�&�&�_���N�|T��`8��Zm��&�K)�Ya�&2�H�z-S�I
Pʎo��L�)�1t��[���F9,Њ��2_̘S5��B�<ҁGji�D���*�1��o�P$��}�;�D���b�����T�GSO�%��ަ�}2�������tXw�7���[�j���e���Re���.~�-�b*gu�:vPX�x���9�>+�G�@��X�7,�"�G"�t�8	W:u��
k�q�^��C�ŷ?����N-�i�/u�K3'a��W���1]ZLv%Y-�h��W2��
������� �
 �����J<��[�r����� �����We�Z�≤������VQ�#H�s�E|�V�b?���Njb���
�(�C�8��%��5@��f�G�~|��b���}�?��'nD�cV�)��Ցyʾ?�E�k����)n�_	��P*y�*�߲�J@)��Z<�[��MAt�	�bڈ�F�3�:	�g��D�A
��9;
oy����䘈W�T�-���Ң��Ǭ���n��g�3�ˑ΁�`@�6�?�����}9E�ʪ��eiv�����YVl�3�~�ߍ���F��W��WH6�!��l�,����ZG���!�����7~�u0Y���c�kG���&��	4`$V�m?���D��!��^��s܆@�p@�
�������`�\A�X���<ЁuEc����r����\=UX{ы�� ?��>���iYl�)瀷�2�6/�:F;,��Pձ������O��[L���_8>hUqQ���>!n�P"��{ɯ9�z�˸1`��0o�;54�@���%����l�]C�4�}��b��!�U�@5R��c]�/6���R&��=���$E��(�B�Av���}֒@�]%�U��~��
-��̶��� �ԥ{����aʕ�=,'С�� d�����{�6��w8u��ێ{Iu���D}��Qm�m[p���)�E�U���vm�C��"5ț�k��I8��?�w���eU;AA'�E]8��n�p�Ql{�D���,��k�IEms����4�seC5�o�+��`�����������kyS<"te�J�s���T���f�-�ɴ�pY�v�b�s՛������>���\q���1OC=�P�%��|�`��~����W�(�w|�OT.S��:���uE�2�s��Y���ꎕJF�)=A�[�F�v�bY{.�?oϤcP�����"+��~�*�j����n"�}�}�!W��5iyR Yv�:P�gF��]��@r�kUi�ڕhe�1�xGJ�c�����W���8�ӥ��xPeA��f��$'S-�����TF����m >�a���t��z�Zz���T�*���-�U�%��$�k�&n��f�^����'�o����謜PV�p�?Fj�R�H�aHé�lQkx`K6��W��'}�e5� ښ��Z�k���.��W!��1X�Nݦ:��?M#�v0nH�o�e���	�qt��-{��sK<�X+mC����c��*�?�\�y%˦�H\Ʋy?�^��fA �ź
�L���?�6R�8� "���]`
l�}��{�9�*�A�y�~���@|ȉ�S[p�}�ݼ��ކmh*e�4�A/�����yȖj�*��^ݳ�rs�#�|�����Z�.��	�%��jcn���'��_�j�4Z�XL�8�Y�(0�����YD7��P=�o�7�tj��F�f�AMR`J�#X����p�(a��E��U#�z�Sih�n�I�ϋ7�R+�n�ѿ
������H�v��o��g�h��7c�1rQ�R\V�U3m�<fF>�*!в�*��QM�1�Ns���Me���U�p���$��`�\�q4[�9��
y$���P�ѝ_���a�w���~}��2�X"�Z�`�����s�w��+���?�A���I;�p�J���XlxVHYEB    cb82    12b0�m�e� L�ǰ@4
�*��jxd���p�[Q�C��rc%JB!�b�����dǪ�>�y�B�(�d!��UC\�xrsLc�E;A�(�)hQ�#�IѾ�Ċ�[��"�KI�d�3y���M���[jK�X^kސ}�ե�;i�{������R�m���-��:�<t[���=.P$��c�æJʱ+I�~:#S�%�:6�O��
�c���_�b3`̔.r���?PV�~z�[*�����)�o�~�q\����G��I ��lѮ��|����fߡW,�d����z]V^L^G�J����"�0;K-���	��%�4K�ad�w�!m/�#��!s� �g��ר@���Y�d�9�/P�gz��%`�"�(09��$b�g�[�������0�n��Y�% � �x|;��hQ�n�G�q,�$��U���kUdX���koK��8�+��5��ɵbfM��Rc�p�|.�¬6�b�k��-��Z���t��G�f0# '�L�h��݉&�w}��\��G����5�.!Q"0���'(��>C�;!d%�E��[m�N��Q�%P$(P{�A/oύm�.���M�_6�mb|��E�%�Z��]�|b�ʈD٤���R�W}���w��7K�ond��C�vb|���9M�^H]"FG���
�`]$��9���[$�P�� B��b&1�XM�r��.%�p�b6h�������z�Ƌ�ҏ ��}Dr�����\���UQ)#��?��j0,RKz���k2!=#hS�dT%
��w
7,�zzvxA��>��A
��v萃Џ~
���G�Y���y�H����9��+:�=^����++��z��>�Y��x�
��6�a��D]��*=U�+qhj��_�U�
v�&��8��#�fһ��RQE��|�J��eN�|��>Y��
t"��%;��������f@~���	ث�	Dt��h�	¹�� ��aqm�Dp�����߬d�2 z�� ,sޭ�]A�v����dP��҄�/�# �h	�m��L;��-^���ŗ�@~,��kz�=�SU���&������e�a�z�X#��#�!�u�W���m���'�O߃'XN_�E��?�3�w<��b($��&c%O�Z?�0��m)��ԭം�/�U$��ޤ�f?�#!��H����©=l�ȃ+�� �
����1oq�����ÖȈ�o9|�>;��е�5���:3�^Nv�W�����4��5�)M5x�/�GI7?-C�=:�ȃ�\�G�a�D4'*���b�8W�"a����F,�J�r-�˜^_�C�a\���g�r���и�"��ȅ�:62����s�I4����.�c�I�hI9�8"Q��J8 ���7 Ý�/&i��6�����y�Dh��Lw�96nǃ�v�sb�#��rl�~�,�_GI���bg|Hh��BV�l$���}������,B��ǭ�4F�(�Qj �m(dMz�I�D�E���XnC��-����U�8!%�"E�`�P���e�eH�?Ȋ�}��#٣zR兞���_���Y�B���tȲ�|Z� Z����T�(�b؜&��u�~K���Y������a���v������nu��Y�w��S�gkb��v�����o@�*����� H�x嗰5��5��[a��GUPQ�����e`��*C6��Q�=ீtě�V�릡%�Zd�Kبʕ*pWt]p�3��H����x=M�̈�"���륓hUS����ud8o�?�[K��K�_^�u2g�s�'��]���5���ӣ7�N��b�䱍�a#�ʨ���x���^�~�U�ɀ�?�m��M�O��@�LF��2� ۫t�]t^É�����Kv������������A�}�D�EH��.��}�����/�{��
^P��*|Q%�+��5Gs�:�����T�4�xN�Qa%V� � {?@��,�
��or2�F
����l���H]�l}U��K������W0U�s��b$����)sw��'���B��_×ծ30��	E萔Yu�l៸~u4{gE��,>����K?(X��OI��|ϊ��$h��w��1����3�8�dM�d!�{Q��7�EJ�I{1�~%]F��/F�+��4��R��-��𙺬%�WكU����"�^L:��Ĕ��l �����|X�5KG�p��a֏G�mZ#��
#���u�-��H`.��c)?�8�R�g�K�Cw��Ѧ��ے�r�i*�m��?�㩧R`f�V1rJ��y�i���2Qr���f��p���Ÿ&�r���tGq9X^f}��_�@Mc8$f�a�'�Z�"$��7�G��^�_U���`lJ�,�~�4��ۅ㍁Z�>H�A�Y��L���6��!�k�9��o�C�~ܝ��C ��0�> �vo�Z���K��{�å�c��R�����C�u˩@0����\s��
��Zy̬c.TQ�`Y�.&WU�iC�Qd��X��"��� �8t�!*�܁|%Uu�h�b��0k�����q�3Vӽ�NK�G����e�������5�
[����"XH8�t����,�A<cɇ�
�#c�.�h%Cr�i ۚ�D�� {m<dp,��9�=��u����Y�FTTQhz��іt����.*��4�2�_�U~1�wS�n(�;�t�����v�8� ���:K��,�-��H��v�K�FG"��{��˭Wa�&t�߀�Ty�^��@ր��O�#�H ������֫%n �C�/������Wj���7Ϡ"� :y�q�/y!��綅1��YR�ҏ�c7Z&�&lj���}TX��ɷӾrW}�<:VY�φE��Y�Ǽ���9�?��oؓ-�
����
�u�kC@Oƭz��/�@��=$?�ZG�����\`�7N�--�2;��̅�����ݤ��d�ymG�>,����J�l�G���9��fѾï�&}���7�����y�ɲ{�;�Y�t(?ڤn��I(Z��_��R��y޹!�R�v�� ꉙ��e��\�1z��$��؇V��0� _Q�t�_3X<Dﶺ�� �b��[��»�bGz��іϕ(��ǣ���xPҲO��S�U�Kʤ~�U��WQ��e檎^=$\O��kp�t��j&]ך����0-�34��uR�ޑ2y"V���
2-!�Qw^���(\c챌ZAR��&A�Ƙ� ��(oAv��%F�٬S������x��=�s#A�����������ԧ�M��3� �©�t`��/#N�����J�t}�$vǿs���pϵd��Ν{�~��W��i(t?d-`����86Z�%�j2�Ty!�~���@���'Dr�(�Y�z���ج��v�;�l꘤h�w�?ש�u^ta�7�/�����>GP�O�[�b1��E�8���d��YC9".��]N��QA
%�_��[��G �Ȗ;�ޑm�����nj���֙k�ͤ.�6�a���7�x�6��L̀�>A�@��z����h���8�;�k�f(�u�]�~t�@v��\nN����X��0B�����ݐ��<_�-F��U��|��5m�8:��m��mpw��}?ٞ���90̵u�YSfG�>��ڰpk�՛�2��5 ���{�a&��/�9.��8��w�8�H&@�(�*����Q�Ri�-g��Ц�M�{��
�%���������<G6RyQ;�gez�H>���24{���G2����0"��3��Zk�%�Ԋ�Ԁ\��K��٫Щ�[v�������u�����/��$9��SֲS�0� ��~�56 T�D12"�!8���3M%�U�V�X�\�:k߮oi�������v���g��4vDH��H���V�IƳ�����X��2qQ�~E��x،O��ޙc�}w	�q}���3���Z��V���DQFȉN�To��76A32s<��@xɁ���Im͈Ӟ����;]Jv��O�bed�wՆ�i���}1�6��I`��㒧��D� 9O��Io��[�� ?��|Y|_�7æ4g�wJh�JB�-�a���!�`J�By[q�u��o_EAN-�@.���m;U�pی~��d��FB_/d}�"�v�)��J]���������Q�웂����X:ҹ ��1֍�Ֆ�cij�[�-�"e� ~�2t���V0.}:�2�ç�s ��Ŵ��Sv�S�i�Wc9�p�u�'V��W���}/��ϝ�@�A
�y̘V����/����e��]�ؘŀ�&��g�Iv@�
�Y���?|��_"�$�LDI��?���[��{���F/ô�3*j�evF�ʳFkK	;{��C�a�`�j�x�����rz�0)��-�$�\b�'���55k��ݿ9�_H��8����W��=��׷TA��Q���UN_��cע}W����d-4�&�𒠚���\��u�s���.~qN8��t�	���|�S���yv^�������>C>r����970���B�Ʌ:�J�TT���v���*������̕`|�Yv����o�	bBҙ����<|��l�Q�ɚ��N`����8�+���;�r��<�[$��y�!Y�Q
��'��x����R�hG\�w�>*2�≿�Ϝ$�ޱO�{G����=�L�>j�4��E���캲,6��YyY��ӌs���1w�y���
�l�$^2"�\���&��v]�z���	yC�,F �rP�`�_BU���z�=��١%��!�6����%+*k�;�|w�