XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���)v�]w���/��p�����٬x��ʢ;����iCkSj���/��|:������l�ԩm	A��e��{�͸��Rs*���ڟu�ˮ^���pR绽� ���Pr08�����:.l�� �=r��CG��~T� sջ�Baih<>����,��������|wy=����8�O�,���" �b�"q�_>�'�_�D��L�R/�����-���:�Į��<�a}�d���jȣ�$�����ΛC�R�L����F.A�]��V	^S���,���l���V���ZMd�4Og��$ �����њma4"��)��`�*�PK��KMR�O6��K��t�c:y@�Y�a���=���P/��%�vu���jc��w���ᆌ�}\�@��Q�����2��tnp�x.f�'Hu�q���0��k�S��X�u�$�)�JK"�<q37��oo���/��a�gm1����l���R!�mױ���sc{U4�@T)O�on޼
������pĎ�T�!;~��j`-Y����(�����e9b��%	B���������rw�\INf� F�?�����n�8�V�)��)#G���ً�vy$S��͸�儞�/��gx��n϶I��E)Z̕W���,ݚn4f�J�V�k��ġ��ZA*�,�J3e��4�L�X.Zfς�A4��'�K���(�rƉ!�|��$�o�*l��j�j��]�;k�r�7�ϫ�u�tv��sՁ&9L��"��1XlxVHYEB    fa00    2560d1������T�QK����i$)��®��{·J��Rq�̂�S_��rk������o�詰��'�����t��ސ��0�c��~��s2R�`�cnF�CS?	z���M����u���vS�� ws@��h�<�ɗ<U<��2UIc�uЖ��9;3���;�m��R;]'�ц'��9�r�|�)�Y�`������Q҃�tt��q�ݓy��-漏��Yт5�
�9��Ս���A�/,A]t�����5�fj��T��V�k=���4HPpa>��5<��C�?&���dh#0N6~)��Cď.٧��G��D���������@dbN���"�+P��ܽV_��շYp�$*�eq��V�H��	'�|�o&�gc06�{iH��~��,(n�	�����R�խ��& �����[.�Ӆ%A�:��J:��H
��l>ۄ����.��4(av���jUfb���1�4i�3�3b�!%xp'�l��F��
H�e������g��	X�D5Y��91�@�,�{S#����[���U��WD� N��OzUĎ���/�;ݝ?�-g�D݄�K+9!��z�ƀR��$<9��H�gt��[� '&����fHU���8|���l+"+<�#��Z�Ջ�e��@�?�����%L�Ύ����������R������s
�J�V$���%�Q�n��\�9�*ol_n�m9H��w���?'�G�=p*L�$sV,?W7�h��X�9�l��SC�J�����0����WN(�v�;��"p���~�v!��ϊ�gwnU;�œ�R�2��EpJof���v�����=<�ş=ǅd�J�U)8�+a�
��r�h̸]�z}W��{Zs�f�7M<�RO��Nz��]��)ͻ�*�v���2)d[�K�Y��RJ�]����h�G	��k�\+-���&�B���*�vR�SИ���=g��w�
[
}���ϰJ��0e+��|�PF�/@՗���N���{�cq � �0̳(�g;s�E�؆b�D
����KV�M�m(�ؑ�]H��7:U�Lg��|X�*�Z͉�g0�f|H���YJZ�wi����b�P�%��˛8!�����=���Q�,Ѿ��DSb�<�s\���7�������6�ug�P�����^4��~��n���7I�-���P��l��:�D�K:���#_�����9�s�W	�踁r,;�Xg_��E7���U�r$>0�G͈����c�%p:�c���PŬ�"�Wܯ�o���.u4��y0�=xk\��7 w�L	׽}<Q5'���-64�7�.��Kf�J����3���Mwϱ\o3
��0���W[�o��\M�+�^�ȸ��r{S�,�N�+RS��ٹ�O�z6P��jO(��YA�Է�I>��
2�[��	�c�V"g�Z�6[� �M*Z=�b�����xq�!��8ey;�r]B�j
�A��g���	H$�)�=N��\D�Zܒ|�����u7�~ݑ���I��C� �א����~�=��0IǸ�/�9�}�-թ��E�9h̛;R�8�mK��MB��ҍ1�n �};�ޞ�d	����-s���z
��δ�7��x)Z�W�bs�񙙜�Q3(����5⽙"��{R�nhh�������>'���S3�ίÀ0����C'��~�%�$P��%u��_�`���_ᶧ��g���J�Q������O����ng6� !���t���6���rz�.8M �Y�$���C���6��-LV?�����'e��'���S�E��d��\�B��y�$���s}������:�H����L5&�83hz$��
*�eD�G��<��QN�+�c`lz2�|��<�����!H���s�9Q�w�z1��$:�[I�=t���s�L��f�r�ݵ������Y�>{���fһ�n�L
���V����R_�<�����Q�&!4� �p1c��IOҦ����իSMd`�K�4�ٮ
���N¾�|;TѶ��˂�$S�K�̌1�����:��8���{?{[&K4��_�y.4b�����̉l��9����\/u������(�Q�L>�F� �\0�]�tV�o�l����<����&�*�9�s߁X��jE�L�A4EH2�b`?Bׁ�+r�>.���@"�O�6��p�HߊgY��BU�N����B�/�'�_�@�$��4a�fS8N�s�`��y�ܟ%���d>{W&��U�V�[�����7 �*I�2�����!�ٶ"�<��|'��S�YA��c�
иy]e�"��ۖ�~���g������c!��:���P�|{��3�>N8�Pej�d�.R�DHv�Ձu��\��_�\��-�+'y���Y��T�6g��!�c��ۂ�v�_�BQ5oD����GIo��1�M��s�$����fF�S<5y�Э-�*`�R�����q��x� ���H�(����=��
��I��:��.e�[&�ʕf��s+T��{LM���k�O&WH�����	p^��(�1�E�1u�W���ZPgz��W*׆;m#jdTXA��~�������6�J),�=��X7��p�7jr��£�ܔ�%���O�
dOv�ɺ�;��R��v�?����!gفZP��~�	�K�s�1?���	���×�� S�Z�U���H���<�,��3�Ql�c�ߑ��tő��wNQX.�����h ��%�֋}�� u�d>B�lu`mȑ�,���}}ĸH��[�����~���	�lkV-�����u���(�k���X'_Bq�3��GS���R�	.���4�Ǣ6���޴��ȩ,��e��PqC������iH3j�N+ۡ-��=W��^�(��{��`�r��o���*��q���t�+X�^j��J�v���4~M�s"I\� 2��"�J�oˇ+��M���L�g�����rf즞�ӛ��ɶ�*Rl��
�G��^�)��ZX	��@Q�������Tf��z���$��-�Ɏ�av���#���+�e}yD������5�	��kٛ f+#<���!K`�1��F�ۤVR�t�qH�qA=��Uןz6e��P�9��7�'��ћm���,/P�.�"ܫ�F=ʼ\N>\q��H�ή�O#� <�[�PE����5�#6�|�]�����`R����+'��+Nݫ�����y��4��a(z�,�j ��l	�Ys���%(&%C�6�.�g�kTI�`��~bU�V�TMS������u�9�l�*k�yg�}q�c�����/b���q���-miUh���R��*X�+�F#Q��� Z��������$�5)���[�3�\=�N��Ǎ$�!/�@Wh�����/��½�R{4��Md�AK��$$�[5	���_���>\f-xw)<U�����E-s\a��Y/�u���ףG3�tC��_���Y*ЁNA�"�Z�x����;P0Գ��{�TX�M�]#rjH�(�!���:*t��9.\=t#���0�.��C*d��x"_vEL
�x�Ǆ�P��K���f��n�/�Fwc�3�b���>�λ%���B>t2�',8�5_�vP)����l']��)�T�<�H�:*$���K1�4.��a@��=�A��� �]��~UD p�n|l�ɰ/L�'NvD&�)����b6K)�À�zCZ������������#���HS)uߑKD�D�m��ڡ����"+a�j7Nh����,����I�'ƃ����E�����q�m�|6�4�Z��0F�h���v�?С�r{:�41� ۩�� �!,BXA!�*�!� ��p9�>�(�H���ysb�l�`�~D��ӝ��6�H�3't!-R�:���&}U�^c^�(h䲈��ƠFO��o��Z;�Њ�ODi:V4���*{'�&1oiP���W�g���'7I�y<b�I�&=Ȱ�	<b^�$�������mɕ!s"���*C����{Qh��qOzW��#Β�R��ZT�_ސ�؋���f��W�Ȥ^Wo�s�3���Y�!*\g�66*��I��O[��?�҈�_a]�*�t6	��K2�R#@Cg��T����A��חV�׬.��)�؞�!���fO٬Z$o}f��i�t�^�S�A���1��@��d��Q�BN��v"� S�l�z���w�j���j8��R9G�7���n%hC���P̮nh����n��	9����0e���9�[������
f4j;���D��ls�'����+��ƚz���Ђ,�$��D&�V�1H�N�Ds���y�e�c�u�1�)/$V
4%wI�L�^*4�� ���u�*:���^�j��l�����`���k�J���>u91����!_�"D��R�?ζ�����Cy5���27u�_n�7�1�*���u�x�Q����A�X��w�YrϪ�%�G��e�m��&�%	��eP[)IE2�}�H�h�b*9�ª2�^�x䊣)Bd_f��5Ia�/���$L�n�4���VY����ဒ+Ƽ-vM
B��ߡL����Zbo&KGo|�Ew��6]H*����.��	�S��k����n���.�m��O�$8e��t���f�&�4������ɓ/-ĳ�0l_xU��*����
�'�CcO̚�D\���z@7A�ڋ�n{�p�F�1��E@� m7[Z����7��4@Y�#ż�&�x
�|g6~b8�.�
AE������w�����}���}w��2N�&�:Gin� �w�}ځVVT�� �=��\���W�q���n�@F�@��Ԗt>�!,/����s�{A6z���I�,i��̀����Q/�g�����Y�+�� �w�;�!+x����~��/�B���_Q�����&�Zw]� ���'d������8�-�&�V�>��C`�����8J�9�Z�s՜��^���p�8`pJn��1f��]����3���i��e7�9-��~X�m��L�W|YƱ*=x�#��?;����EyT��"f�e����`�.�6��H�t<=b�W���>ڶ$f�ԅ��J1Vug�-�_��؄�%'��ЃY�<��;��@�d,�Sz��� �}������T���
�J��S�8����3��j5���[���O��	�+Z�(����IpX
ß���� �պ���E��,��ˀ��G�������/^��� ��cY�(�-�
b:��x���/)�Q��!�/9��	FXv|���ܠI�4��F(L���*N�Q�c��lIIFZ
[r���2����f�>�x̵�N�C1��D�� K��
ْ��CsD�M��#(2�0o�S�����i~���l��F���Px"�#���YUD*���N�E����Y
���G w�HEϡ4r]%R$��&
S8B�h_.�R���<Ψ?_8e�Nx���G�����1�p���������l!R����/}��V�ӗW�DN,14i��h�y	���ǰ驃Tާ������<7�Q�P���g�hή|�U�6C«J��E�ZÅf���_�[Y?:萤�ft�{X�M$*?�l���ʛ�J*�	M�����*�����7`�&�;#�<u�'2>����"F���HqX����(A�r�V-[|V6(���q� \�lI�?~M���t�ɇR[ܠ�]�?�rݐt�7���Qyu������\�z�n�P�"!�ᇄj�G�|��WiM�|W�6�/���P��;��h��}�����>�ʦ !�6��V�N�֗v�Y��KL�����{t����sy�XҮJ]�V��¦�.Q_�M��+]�d�\�H��=���$1&����y}ꯤC�EU�'8Z���O�a�H��8}{q^jk�JSmO�y���/�8��S��v;F:�V��e`���X#�bZ�Ø\�rG�*o��w��C�M�R}J�!#�LHS����h�<ǻ7����Жw��{u���R*����{�]�����T��yf ���݆O�t�����������Q^@]w>�W�)
|<��٣C���#�	X��,��48����u5�L�q2'ΛWdMU�\�V46�8uKm�4��U)Ӄ�h Ҵ��z���v�Y���#B&x�<,Ǉ��\�kJ��1"G�"x�����g?��O�t�.�ca`�����ԡ]�)�,F�n�(�T��fg�m�TsTz������vƋɥ�M��7X�Ő��`��A��a���A�F�F7s>A�v�,ԉ[�a� ˳8=�n x�����|7y;��Dh��Qviw�z_͆���E����o���v!>UK�0@����(~ZL�%���D�ֶ�����QҸ#�$�#tW�b���$�,�2	� �Z��ǋ�EL�Q0��p��7Un&��o�s��j˩Pņ&\E�����1�|Sg��J�-�e���I���c!��X��$��}�"Lh.�����C�1�����Ov~ͱ�ğ ���"rA�,��7�D��\E^ ��?'k���y�m3�Lm2�6�L�Gy���`��A5k��H���يi�E�f��aR�k;��y���"�a[E��P�C>�~�~y37IU)���j<>l6�1�=T�\r�V�=��w�6/Q
�o\��u,��.�$R���ٖK��w�k�K�`�\����M�/e�r��^.Lr�3��Q)ٌ�哙�]*ݨ#�]�W�$P�jR��;"v��{�e:'����L�����[i�|x�7K2�l��IT�����e�����+�Ɍ����*gmnFt�%`�l�������)gT��=�X��v���f�V\�*���h��[Ҥr)��F���B>y�D�Ӏ%���w��{�RL�ɲ���2��7��mc�$�/a�8d��@AWr (ݸɔj�`7A	��E��oR8ź^^�`� ��N��}!�����e�����ds��E���*�53�ec):��ecj`^���fe�����8{4��-7pSg+_bkD�&G-*6F����`�U��7����V����b��2���@l�e��b������ɹ^A��+Ð�P�m�ٗ\���d��1���y�˷�%f+��ZH�a~AU�;�����8����W�����5j������N@Ǧ��2O#(�FJ�s��������K�:s��� /�|�#�(&8�,��|��Vo�}�N�a��K��T��
����@��O�C���!�j_��k7��@V��$�Ј�;g�)���V���������_�X�G7�otݣK��q�����@Qs�zAp)g���c̆w߲��<ט����^��U7`e�H�S�w�T�~�X�'��=��h���}���SK��T;��R��������Y=di�ast�mG��f�ˣ}^��H��r�+0�s�_Ih��v錼&�A�C���3x<g/i�*�ψǑ��%��t�`�@�����	�Ӝ�Q��t�'�����4(�갥e	LԹ��T��yi�B��Q�>�P�3��*�:��V<qަb�0�N��K�����#&%X9�ϥ�0<�6�0�m GTXm!��Z�˲�6�(,Uߊie���
[/�����
�Thb�J� ��[`��!���&�K ��~y���D��7�G6H�=�+�������#;��b�Wׁ$��f��g��<��W�����Ln-���x����AȨ�c���9\�)�����d9�,���5�'�K���3L77�K�4�9�`[/�F.+O�T�e�a�~�	[���&����%��!�m�L�G��$9��.onґ�����n�l;U�|�o��(���1c�@����ۥ
S�.x�� &���!�V��Xô\�Ŋ!����������1[{6�*�ğ�(�4&�D���鏴:�r��b��Ͳ$]��W���<�r'����ov�����7;�41��d���I���:ic6��!!)S<��A	-}�~�r���RZ#�/���Y݊&�V�`1�2�B����w�+Ay�?�iku�$ɔ8gV!zAz��5V����S�=���؞���S��1JX]��"�Sӑ�VvWb��z%�{�=;�:JB��\2��)�(ӏ����ǹ�/�]�bAw���Ɗk�w׆U?�S=�d�����=��Lk�1	
�o�k79rG�l��)�P�>$��<�)�ҭ�Q���;����D�_��}�x�O�r�ھ�%"�sDOu��s��H���=��XS�9l��T����J��2K2{�ظB����@>Q��s��eV���
�,�:�P�R�tUt��_:k����SEK�����#���P�@P<�A�('��Aݖa�I����^Tfs�F���G���O{����穊������M�a�8���{��وN�3��Z"�a���s��?^<�܁%x6�����T�a���s'���D�CzQ�0gC�sQ&S�q!�`Ԣ�1���n��ɇ\in�~�2͉�%���)�O4'��\��g���bwVE:[e�7��C��k:�P�(t"�S�rfY��Q޽uO�-���������nw߀�mP;��x�!�N6��wj̎6Р���ޭH�{��l.��X��z�J�����s�ɼ�C1�Aa:b�����~���L���' <�j�EK
le�~;���
ʬ;�f��1IV�Z�l
�m�?�ƃO�����k��.k�Y\����0�|����wёj�{��Ɋ�)���������᱀��O%��`g��ʏ�3`�JIO�M�J�z(3S�,����%P�4��
���rB�g:8$|Y�HF$��u��Q�?/�_I1K��X��f��[�(������bDVZ���&��/���£E�7^�����5Ƅ_��Љ��}>� �+m�.o�@� �/��y�E��й�B�yq��;�B�b�/D �/����R�t:U�΂L��t��Q��%*ѥ��A Q�7���V���R?E�g�W
�ܳ����]!�re�Q�ꦮ%�p�Gĕ��s	��EEfN_����c��j+�����zYu�Ӯ�K�U~��l��h�a��V�B7q�	-9ޏ�bu�?�	�������V����q/;u��҉��j�*%���O�ƺCQD���W0x��*��Y_��e�O/[P�YɃ�G>p��4��t����Ȏ
��|��Kt@�n���`��'����Xwn"��"|;�[v��u�ܫ�ե�o�۩��O�F�`�a\d�"(�s���mڠ�ɂ>��<��%ۍ���=�7b���=�舌%��ۓޱS,J>]��j�6�ى�8�Gʒ�Q��U%m��)=��iM�C�qN5~��~��nL��o��g3Զ��9����>XlxVHYEB    fa00    14b05#��
�/�>T:?!eZL��V�*��g��Yj�;6uT��b�g��/"�������&6�c�ncҠ��d����*&�P`+`�￟�%)�2%,�9S����,�_&�6����w����C��sCx�4{���;��� h
!���ֈǻ�Yiu�&��_Y=!�9��Cy.$��N~���>r��0J��)��U��3����v�?�_�;��n�񨪂3Jܝg\��ʓ�K���r��j��,���D�r�<p�@�ľ��@�D�h�� �����������%8��+CeȲ�m:8ST�vt��#K��0�~�$~�g� z�H�w���mR�"h��܀cg5b $c����>"�̪�U|���Ld"� �d��Ļ8u�Fߤ'�!(�P�hϖ�!���n=̉s�I� ل�N#�G�X.�����cfKq���o.θ�o������CtV���E�R�3�A�$0?�j@-��G�ۀ�Si^G.�o���t��M�cn�z�)5�������f�B���o㿯3ع��/5Z��I��8��j�v��9kwѠ܌v[�@;�zOf�2�[��λGSYv��\��ɤ.l�lݷ�]�Y����t��Y���r�&��T��'�F���GW����ڀ@t�uI,P�3�����8��d �#)6J��r|��bo��R�=u��R[�\^&���|6�-Ìj��x����&d�T6m7�i�P��~X�v)tH�0��!�1u���nю1�*( :U�0Ĕ�Ė�tU�S�$�}J�`%��1�5
�������TJ�g�����^�K�p/d���U���zw"~�_�OI^0����S�@�Nnoj�c��+�q�WU�zv����\Lb�PH�(���F����>�����d،���S@�$��Z]�+6G�{�פQ��}B���j��Ҷ9���J:�E�i�uM�᫡q�u�LsƎ�mb�NɾNe,F�<~#�o)Ǿa3���T"Ok�)t,W�V"9�Y;-��ń���.�۩9*�58TZ|�.Q�0���[}�8���X�E0�Z��Ҽ���q��ݨ��&25(��n&��]��^+��Җف
?�Um'�������=���W�w���^U4�\i�<^�c ��-a�y:y�m����jl�(n}�������(h�����C�?�)��p,��Ŭ��%�|{�K+K�� �Q3�B�����l�'�:��5]Q�����t\�@CO��s�SM7��v�8w��Rf5I��Z�-<y&�o�0]�W�a\��\>[iRaT�ՙ��I�:حO<"m���l��j�Oo�+�OwZ>��qJq�'=��C4T�'������IߟlE�t�^���(@��Ac4X؄�̘��=Cy���Q�	�.94��{�)d�+4���D��(r�d��Ж(�quh�B����<�y[܂\���.>�;���'��S䃲;A�U}���{ȲjW�^�^��3�h��D�.�����S{��!Ӷ/�.�C�Z���iaP3f�܎:�����4�HE�'�/uz����<C!�7�\���<-@����Y
��/�c�8,�_�FM��N��Q$�V|h��<rT?ք�ď�J�j?h��(γAq�Q���Rc�����Z9�M��=��z�G@y���`1$�ru\��UYҙ$�\�VKϽ�]	��[�8���]Eg��a�7$T���Jŵ��aE$�o��]�.�:��k�FĔ�В�$,��^�93.�:�L��>�wi��F=2|V'�	UL�[��y�bGliG�v�T�a�Ulq~Z�ܳ��R����e0�q�U��ү�謁V�v(��=�R�V�uw[E#�`�}a��4��B�F�%����L�P�T���p�='��Z���n�<6��=R�h�zoa�`qx�V�v��o
czB�^P1��4B�f�Ƌ�;����,�c���� �� ��*�­�$����AbF�����?��56h�Z9��Ī�?m�ɔQ���8��欍�
"����t/����P�v zЦ�b?�ߤ3�W�c�l����Ic^�Z�Ű�VG(�E(7����r�9ծ�|�b��'~���ٌ<~�7��F���ߓnNc�<1�Z-���,����e`K�2��W~z�a��T85�o�H��z=L�C��r����ת|�M�v��K��}�~����18+�%E��Nd���_�H�hj]0da��F�;��þ�l��`�e��7W��R����3�c_5���e�dK����ϡ@9M%& r�3����$]��$�@Z1�2ș�<uLjk�P,/��
��}s��؂m� }q}	�>Q�GCE����D11T~�'��^��<����N��"���"����bҌqB1�c���^V8�H�9�C?u����[�4�ֿ�	��{�ap�	�;*͐���q��?�0��8�ЩВkKR�6[j@
�%� T�rA�~\�Od�����!�D�J��j� �p �I�hi��1'�D��])
N��r)?z_.���x^s�<ԅt~��'W���9���E��U_I�Hrd�����6rs>�9!�g�Kv���[��bv��+:���ʵ�{���]ss+=�` r`�u>��ȐPʌx��xm�*#�n��縋]Rvt���� �1�ȧK+�%��T��ǁ���>!��:�� �����ǪN��~�����X���k4�����R���	�ލF���oa7#��_�]j��R�F�TZ�ښH��PZKM���(��**j"�x�����v�'�#��������@/���[59����ȡ�s���稷�)({�k� YRV���)`��KP����Q��h�X@�Q@���A���؏�LZ�����7��{fD
?��G�J������1��M�;B��|����o�̏�h���W-��'lh16��Ϭ*CX7W�@�d�1� ֒�3k�O���uU��^��b�b䧈�XtgZ�:��%�z|
�]фX�d�0x�����C�i��$ŉ�zs�}Ab�j��K�n ɫ�P�\�8�a�Ƒ�y� C��x{
��F�K6�����s�����USd?�3Q�5��}�|:2�67����$�17��� `J�h��$O�]����`��N�F�v�_����\q�N	��#d��$%0!'���)X��J��m��W�^ �9q&�b�ؒ�6�d��_)L�&9&�k�V�o��U�ʴ$yŐ�y��{ׅz�+���'4t���8�.%	.�}�=�c
�'���`N�e�H�$��(E��W���cG}�4���FǛ͘�'�ch*0���#��L����)�h���ge?[	���9� �O)��P�i�����+}�h����щ9��0�ɥ�:Yl�s����JR�\�q�d8�sD܇N�lR����4�st�ʻr����k���oW�V��	�z@E6��X��v�N���`�������(�:����:H�ݍ鰐!��������:�	�Z�qC�d���Qj3.�$��{L;fRf�u'����LH� �V  ԋl�	�!�2��ʩd)8��r�	T�ӡ��Y�0�WwQ1���UL������������v�1��&��y�\�Wrk]M�Ļ������4�������8 �q�]vD����[����[�w�8Y�2hw�Z�U�U�oEr��0�w�P���sGf��U��
\���1��%C��t���K=��J��=<�ɸ����W�����?;���n��Wq�k�9G?��ͽ�ү�^�$�tXa}�Nu����GO]�mы�� � ��f�1-��M�v}>��h��C)��dߴ��t��Ftw���.2��덑���xPE\���}�￀�A�H<O�����eAw) 0Z���w�N�e/+&2S=i~U�l<8��׍����ĵ6��s%P�L�I°܆�_ZF�Иy�����5鿷��� �n��VLӂ̄G/����ǘof�W��pgKO$^���P��"D��0lۋUx�^&#W(��5�����6l�N�iP%2���Π����)� /�"��;"X���V�C)
�EJ�\̇� Y����.�g"Jj�U(�q]�@��������ų��g�Mb9�E��M%�[3��Ի��cM��+���u��0�qq�і�VŒ� W6R�>P�-}�c��T{�Ӂ߃��|��|�{��y!u1�
^���w��v�̎��}���_�~A�+��ꋃ���͛�jzLb��Y(:�O�5�qM��v���1!���b��l��+��[���YX�Q��\&~VVN����{.p���=�n�f�[�4��P�Tw���b�4�����I7z����?��pJ�=�1g�x�`��	W�`4�4�4��x���(v�����b'�{E����#Q0�й���aF�\���j�*�nF��Q���l3��h�]�<�i;s^dc�[:�ax���E�8����yvT�z3�)�YI�&�Y
F�5�_�Ŵ�8�G��=���/ꌢ������[��ed��[G���d��>�o��C�$h�z��Ф��&P�y�c��I�g�6�cE��arw�X[�+['Rnr��e�y�A���?mѰ0�%���ٲ�sT�a��v}����e5u7;�"�~�mN�KQ��Y���YbΛ�X���}=�&�yM�,��	E�����\/��s�����Y����&���f|)k�Mʚ�<�a�\�9m�a�����*Wl��4�� �(g��*8>�
b�`_{EB�d)��ZּG�Ԋ)�p�$�AFѦ�Y!��(>{L��T�GM�(@��bg�.W���E1ѷ���������{�Fո��SM��A�-�w�ߪ1�$�[NO���U�/R8XV��N�����J�P(C�yO��2�v�,'��W����r5S���o�3ݲ �A)������C��n������WL����j��R�,�aوu��]nȉ>�!n�-��ܭ�y!���U�s�f���Y\G�^ۧ�����v鿿a�Aj)�UI&����?�	gY�M5�y�+Ń�@��J�X4����p\�T笨�S��ڇ�)<�b}'x�N��h���
�B�ߊC�(����J�����O�?TB�M��;Ë�T� 1T�}���Z�����^4e�D5\,`aC�Zpn���$
�4�DI�w?�]�H�_��k�[��k��G�e� DS�߮�����h��XlxVHYEB    fa00    1880� X���{�T�v���%+ۊ���UDyH��Xw�L�͏f�2���K��5��i}�<�qZ�Ɖv���]A�%8�I3�7�wsP|3p��3]9�x��)�������9�
^�˚�:s�Ї	�u �w���>�L7S!N�+�O+Ƃ�fYR�|����v�ǟu8��k��Ak�0�v�	�c��*��#i�d�%{��$2{=x��=�,���u��FGܸ�5º���q�}��"�T�=ܫ�!�wG�<)xM�����hW�8O���M��u�_�D��$��U�M��� 5����PBpE��2p;5M�g=e��	?Sl	�%�Ђ�C��*�rɟ�t��#���� �e��]���g��p����[���
���sY#�����Uя{>}1ZQ��:�ݡ�v	K�4�f-���ާg;w�S��V����}�gs��ݬC�HmUѹz֎�MM�V��J�n����J>�K�9�;�h�1�ॹ�Wga\�5ّ˵��v
~xh�??����p�nt�O��[� S����OF���cEP��(�� �Bd�- ڥ���%#�+�%EF���������A>#�6y9$i]�6�-Rk:�e+����K�s����3��4c/9�g����{]P��e��ՂB�4E�{lێH"�)����92���Ojj�j ����mGa���@�'��y�O�8֌�]�Z0���d	���6[RRA�����x!�6���Ӳ�L��G�����~FL�խ]�sS��I``2�zͶRg��z���[�e} ��#���r���OG����b%,���S�R4��+Kf�$Ц��5�()ٰ�Ç��Z�RBl���+~:�'Up�<�5,����O��\�A�L��0�Z&򸪒��C4��-����j�����a�x�����!��9\R�Sq�˛q��ƿ@�@m?ܨ�� ��C�j�'�[B͂�hӃ�t�Ô�ߖ<��ׄڥ=�C�B�n33��CĀ�O�u�x'�� �s������t�%�*/�$$m�������Y�G���F����f���֯��:�%%7��
��_�Q�>Z�1��G����F���֒Q����-j'�O�(�V:l�*"@EnG���zt��(ELT��gV�>�ܨ�[x�2A(��� Z���4��o�񡻶41`_p+�?SA��.\a�0D�z��	^�Ä�x5�&�
�u�8�EDY�h��/o�:Ss�aM!Y4|�Ώ������������6r�vB�|0=2ql��Y�^BV(��+�Q7��0J����˛�6]���8z���H^.�e�Wh��	m���^��{��\9���፦ӿȟ��K۹I\��N*���kL�:'hg7���^a�2���6��	�Y���Rq���9�=or�����B��`,8����Iյ���sS�l�x��8��Ȼ̌���9�F�[��*����j��N~�`�F�� QG�`�s��o�����S5l����8����y�|�+��6�kz���@�2$��Mt��&fI�BH�����s!X��$NCWj!��:m��L�Z���y�,�i���N]o.h��>��@��(S�b4�	E���
�I��0[�@'#h�n��v5	XU�t:�!A�]gP�Cq5�T1�a����)yLu�P&3a'�5��R�=h�u�뺏KO�K��h�>v+�^��Т[6,;�GSaM�g<V��0Q�Q�9!�<X��-���:����tiN(d(:��`Sj�-�0��ں�P�Ԡ�i{]�{z��SR��rX��VFU���h;c��N�sbrs��N;�D0�xK6���#�%K��()!��Ƶ��KaU �y�3|�S�0�Ř6_��cN��{�q[��1X'=s&�j����E���s����Yw���l>���]!e�S�������$�|����#�
�L��dg��r@�,b�a,��aɇ�6R~_�b�����4I})��+势{���["�.��7^�m(n<�J��D��!����AO�]>| �����,��cK��Y ��G�������꫞Hr$�{�?s�'����Sx�{I&�n�e�;gpM�2��a)��bC�k�A�z�p�왳p�تӻ��'���mXDTW�!�Ej�Ub��``8̭�"B�ߘ�0���&j1s��F,>���ƀ�� :����v1E��ں^������c��]Iz)[*3�6o��&��'�Ǉ�Y`�8N����Z��@t�c{��w9�OJ�D��CƂkLưx�B �5\7�Fi�P��2Ȥ�'C�6@�j$���Pt�����"��JG��E肇��������獳�����$`���E,���Rt��q�}Kv���JM�ч�]7��>p�;S���<����6���$A�B�~�(U�G�r�Q�n2wz|�	���� \��b�����bM|A�7B�T��Bc[���HT	�렑�\�Bo��=]�#4�l���2��	輱oh��\��A[��>���v��p������0�>+6�1xY(��m&r ``����w��3^�h#ҫ�����4+����҂y��`F�#�Ԯ�Q僦�֔�iB�(��r���k��R�����}['w�C掄�yS�}�3T��s}��.���Xy+jiG�1�����݉��kg�;˩Gd�_�!\|�s�ޗ�PeT�D"�.I�q�������LV
�LA��u�/�ϼ����AU~s��s�HB�%�"r��څ��x;@u����&��x͕��Ĵ]�=��8̨��#XI;��e"�.�}L��X}�+氵��Ky��t�ҫ�:��GKұ[���8�kN�1̒�A���md^�`G����;��0��!��GV���0Zڸ\z��6�:%�neM��%Xh R���R%��*_$ˢ�[������Jm��I>u�d�_&��(�9J��+͗�&���g=j}{��t��x|	U��1��oآ~#fI���j���a�	=�rX	�1�N�C p$ݗ��P?��0��6��ߚb��kr����������ZΗ��)�T2�x�^�0I��S斄᱁�qq��o(�Շ�슉�^���M
����c��g��	̸`�Q��	�7�P�d�v��3"#o�ˇAi[@t�3��]�K�/ �Ⱦh�`l�_qbW�Ġ+VQ�>5���{bZ2���I�VK���4K������'Z:��1�K�n�0�$dm�d�+�T:�p����s�*�v����1UyA��I�j���	w�2������
��OO� ��O�8��]��r��L2��f ��Z��`�&M��n�W2LW��7�MwT��x��Y�;g�����Ý3Q8���a^ �`l�YY,�Ka��G�fgݱ�\�Ͽ2��[�Z��sw��F}�"�˦9����zeg��׈D�[��k[s�J���D�N _���O�[x�����~["���G��uɢ�� ��3Tb�i��(�.�O*L�;xD�\߃z�6�$;w��|`�]ڬ:�ݵV�18��1u������|T�f��bÉm�u��օ����ŀ�]��EOm ��t�^:#��Q|�;>���Њ��0k"JbxC�[uպG�:{l�eQ%1�@$��z���͐C@���H��$P�*��x�/G-@�ٱ}�!�oӸ5�=~H��.Gjp�h�C�
�:Gv�?I��e��	�����~e��U��ZJ�������qj��g��JOq�d�4>�C����-�j�O܏��_cGhi�s`�~�h�{&��q�j���f74�>�W��cI}��Pwk������O�q� 
T�@�MP�5CD��׾�I ;����;����Ob�.T��^� ڄ��{�� �%�S�'S�c@�,�r�� �.� X�⿅<���1y���mK�}^��M��>�c���3y�;�d��@�Qx���a�y%]���!����_��W�UbY}a<��W~(l�>��u�3����-k���.Ӳ�k�j(�ױm{+Z��r�v}���*�%���'�*��oJ,�\m��^��~��óI��a/T��|r�R,f��2�l[�](���F�k9��ݫ���jN�+uѲ+ʁ�_Ssnv�O� � a�7E�5?\@��S�F7�Cm��}Q�w��j '�����.��0��YO|a(9�šh����θ�Tg�ی�#��C��/�@|���ފ�uv�+񣒊�um�p
ঃi�'CYt+�{��"[ma[�(�H��,�M�Ou���#�Ɛq7�� �(@�oq�N��+���=>�׉]��z�-s��%���2���#vi���7�kw�l�="�r1 E�,�å]�;��f����2���J�{O�:[�g10[^N�H��lnN��VQ"�7}���Ҏ�B��sը&�wu��6ߍue�E���yCQjP��!�� ~�$a�ªܿ��xɻ�Z���MI*7`�d���M��6��FnZ�lb\ڙwݚ?���*4��Ϭ�e>n��.���' ��τy�8 L{����X3e�AL��JcK��u�C��jw��b��wP�`����wbG�b���2��E�����
����]P.�L���'�Ǖ���]Q��X��\����׌EN�/�^>�j{�W�
N~������Ћ3��J@��TeQ���r[���_ZH�����C��7�f��N7E��̫M�H�_��f]O23��2���Ĉ B�
�Eb Q�||�E��[�.{�1�tWݭ�濅v�v��:��I���@A�3��1�:�U,'=�C���<���Q�7Ǳ����O��h��=���\ɣÈ_��%���Fg����I��s�ԗvh�w��7[��m�2�h5����w��:�P2�>dv',�O��p�����u�*�%q�L���=3�{��<���ؗ��� �����U�3a�"Ln�u<4n�U1��;>L�8=�:�����P���H���OxS���CPdc9��0��"M�����feFf�`��-�)7��KTN���
��:g���#o9���P���F�+3��Z���IL��Xt4g�b�˝�]]ڸ�4�/��}�H-]�����bVy=$�����F�Gn�eEC���V��]YDu�}�+;oH��^��p8��@�����!�۸��E
�]&QlE6%�)ZV���߸���æ�Ƀ���W��mr�ߕ�&�����ͬ��@q�d�u'b���/�U{�Y�z����hS��	%�&��Y�#��n,�s"�X�~cv5`�Kp��t���- ��cѻE�5�I�[��6��G�Q)�X6�U[�g����zB��_yK�`�G� G�\�މ+x�5�Cn`����:$��x=r+�1��΅��ƚ�k��0,�X�:k�#?�c�Y�(R�-�5�^��&���?&��2�[mjt�:!%��Qg���&n�x.� �j�!�$��3 ���İ/;��
� .o�
���c�-"r�H��V%'~3��;���X�#
MV�.z��h�M+t:�]�N����L��z)UV�&=8=s�M70~���C %�⧲�(����&��c��_\8Ď�˵k���%*绤{�I{&�y����@�~&��à'�27������48���a�=S*���9%x�1n��+��5�Gm^}�N]����cȥ�j|=���_�0{=�6o�d�3��������KDdDy�m
��I{G��o��=F-�Y7���rr�e�jg,K�B�Oe��fu�Ë���ټ�g��?E��S���wx1V�mFh ����mDK� � y�ɂ )�;�(5a4GD���,r�g��l��[=�ŗd�W����v��2��L+�>��οͯc��{��{�x�d}�h߻	�v��]��U��G�̠𭷜gjk��9�j;g��x�� �	���JJ��W�H���:aJ� PQ!���
�(mo62]B���,e� �V,��5+�Nǃ�vލ�am��`I���E�6B <eS��D��t�a/�z}u��<�������x���R??�/��(��zU�]:�Fh4�.��c����O}�	����������G?��蠲��/�g0�|T��.0STY"|��A�=�a��A���O��'H�P�V1]����-��
$NXlxVHYEB    fa00    19105(~]�ʧ'�-�b�;Tk��qvt��L���M���D�ً��x�ۢ�&1�� .�V�W9�ع���±�����A���9*��{����?�떁)����$\�#�p/������m�!�k�;�-Hro;���7�����Q(2��J��p�Шi]�scg]χh��

��g�-���� k*l�Y�b�r�9
r x'̎`�ݩ%#+�G��,S�9fo���C�[W���V�ӏ�P��� >���:=�Vi�!��an�xͯ9�:�������z�~��QaW���"���N��%�H��+m���h�r�B�Z���/���	��sjr0Q���5=�a����m���'C4p�D�Ř�v�<׀+��7�<ؼJF3�-ů�� �D|��Мy�мv}�K�}�π|��Zn�[��-��6���vg��X� CQ��Hu�:S�:�=e���F��T^���C��u�\����[���i��y�/�F���C w<�: ���-=��7�
���"\Ơ��3�n_\?���$��~X�Ū���r���+� ��� %3D�:�ª]b��`�
��(aA�O/�@��.�yFtc>l���ʆ�e�zC�C��X���XVL(�s�D*Z�1�}�+���ޔ�#�Αg��7���;NP����f$��?����^@w�,0��N?��n�,�
��uQm�F��o���ފO�D�F𠴂�|��A��j�m?�7c�H3f9{C+I~��p�����V�m�z��v�p���3��f%���=_��	N/a��>�Q��w�|�4@ #�،��0����H8�TW���գ�xz���ʌ.�E���zM�Jҙ�9��Ֆ�+����NT����Nʟ�D�]��үh�Ǒ$@`��JM�0RW� ��Ț�Ls]�tGΣ�k�ޡ:�<
5ilN���VR�+	)�����z
�]uQ(�� k?�:�A�R�D+��\X��k����O�:���ۦU�%EYp�!��`��nUǬz{@�60,/�;��P������+�A��i=%,i)���q�K�gZ�6l�F�3{�2P�_\ҝ�"��u���X�-���QcSv^���
,L�9K�p�^@B���C��sE�,Zq�寢T�YFM�l7Ftp��3�%h�7{��(�΂�{K �;�|�����v�||(�O�W�< �����˪�M�٥E)�S~�=�
���̱ja%�OEK��[����`�sI%�Ri�T����oiAVxٞ�e��j��S/sc|h�_m��;�
�����t|�<�+�z���'��¡H)ҙ��e��x{/X&�)K
{���f��J��5Q��ߍR��L�-w^�kyZ;Nz�O3&:���IL�7bY_`�%f�G�������
.�r1�J�	����?�$�>�tr�ZG�b�p~��Bj�Gz��&Ҥ(%��&$�`��3G���h��A+V�^{c���`U�S� C�hHv��]���'�:�[����Qơ$�-T.\};�#Z�
�<�UU������(޴~�\��ǿՄZ �ʪ��m�O.j��>&Bb��&���C�gF߰�Q�灁�q`UiY���_��IK�BD`�V�au*@?>�����M�d��(1�-dl���^@Ho��=�̀ʛ��nA�p���ԧO�&UXs�M/k��%�J���P�>e�4S�6M������%Ư��>R�]��+����wr!�vCh����|��cZ޳��Ї�(k���-��h灵�U�8_GA��Q��lF����
�R�,�F�)
��n���R6�&�EÃ�8���J���NV�[q���a�V�"��)�u+������g8���YK�D��>��b
?�Bڏ����c������G���R(����JKHP�V��1�d�zfX`�h��c�����Z�G'N����n+������TBBަ���uo��1�4^Y4N�=�����{�_�F(�0%Yy���f��53U�Ե�j'�_�d��(P�������\��ޚ� �J�nÄU���g�g�\�~���~�+���F7���"�)[�'E��=��{㫉���V���t�/9Έ�2��>�0�M�ѹ3��%�N�6K>"��:,_Ŋ�����xEN��"es�먽V�[Is��t�Gc�t\ɏ@�����o=}���	��&z��\���[b��z�A|��D�>���$>6s:L,Pi8�]"��=�.�d�f�Y^����g��F�]g�������
��nK=g�}\���L%���?k�t߼�d�ժ]W�t�l��!���A��e\������L��Wߴ	��[b}���t#��*���s��!�ޚ}��E���@�7��%�L�$��.�֩�8&��)m���A���	�	j��Y��_n't�8�ܘ�"ϖ�#�_^�0i�'�X	�Ͼ�vF.�ރ���5���XV�]���ъ�����A�/��Zm�̼�< [�a���*O����^l)�����G�Doi���E	&����Pu����A�����$q�C�Α��߽�b��@���E%-���̍���h���av�q	,��������?���������o�����јA����$�Y�},f^(2\�\�fJf��Y��9$�B��U�@Ql��m���)	Q-_��.���!���\���S�e	BP[P8�j����Y0l'��4�B�;ʩ�\����h�-o����_�Q��ɼ�~e���I(3�O���5	�`���	^�[(! =���KA�i�}��ڄ�0�T�SQ%�������!ȇ��y9�����N�B��s'��8�X��Q9ڜ�yL@o����o:��s�K�`Ɍ�<���3����\��
��$��0)��FEC��sfC���1ҰQ�����'�j��K���h��p�[�_��v��^P(�&�N>���J)������ܠC�{�l�R���H}�U�/%�[L�+�}�N�3�$�{.��R-_�17kȒf�fjy21<��
���ye������tE0%�k+P�g��� M�{�[`P��1eO�7��u�"+E�$'������7Wx�p��'��hˈ���%��c`�E�!�¹nN1aM�jʵ�V!�B���&䅸����"��P	�Ho��*_�7��N�����.
&��qя%%��Z��K7}L:k�.�������V��h���hk��KO��r�.,^j#$��\Up���@�����|��Q�ƾ>���8�JӲ|�Mr�{��7p��Z��y�ǃ5��T�,zCd���f����3�=��1JUi^��e�p<��W�(qD������w��0��Y�f2��y�P����"8�������'�V�&-w���]��<�t���|�t� ��Z0~j$����� l7��/��]�� [��cw���#��[\�~(��%�I̗�Oحe�Ŭ�3#���LV<1*q`I�U&�Rʨ�PR�w%DO_�����"����9-u�� ����"4x��u:/���l.�m��E�GTj�
y̾��$��#�ww��_��92C��)(�
������č\ơ�]�f���Q�5�h	\.�Gv�QYZ,��#Z]��\���^�6��mq����TX�D�͔�H�W�&aUTV���f��h.0�V����,��̠����6*^��_�]�	���{�&�ݡf�n c�|	�
�6�V*>s�x��C��u#H�AI�h����4;$Uy��,���b���#"x�*�'Qt�l��9�ZHʅ�����q�k]bJHH�/%����b�&\�0���Frg$�+ V��zUXW%�AI������U͑(:$ESs�6J�����J8���\� (Yk���z�%9�;8�>KQJ��I�?��ǭH�  wF���Am���F��fW�����qh稨�O+��L�I|�I"8�J�\J�I��trR�m^�*�ى����8i�s�F�H�e~���8�����A����Y*����7Ե�"���u���-gS�E��@���XjT�o�A�¸o�vT�u�5���?�x��Yn�K����l"��>@�!>�ѩs��}9��8���#1{�}�r���[_��E#���?���#~��(hW�bOj�_/����[���%�����`)t��!oco��}g�R�2��*CUه.*kg���@��P�ZNV���
�hpL����K{�wx*��w�,�po�i�j �j9C`��"����hN�c5�Z���j����fz��K��V�e�=u�W �t��_-��	�~��HZ����Z�1�PO��qZ��L� i���%�_Vk˼ ��؅�M}���HX�ʠ�'�V@V	���H�A��7��Ne�?CDﰭ� �if��D,��k��/_�8�0�.[�ƽp_�����
���HH�snHj�̹2�E��2�yE}�����ق���Q+	�}� 0�%H��Bv�9/��z��,b�<��S����	ʅ�\|eYBf^w3�E O��%g�զT������X5�H��0
����w�h$�Dʓ�����p,]ע���X�\z��_��V�rT�~��(��z�Ih@��V��@:c�"��v���ȥ`	�7�1��u�s��`ʱ⑿P��	��5�OQ߽�m�k��@���.���~e�t@G�V��f��=� �ݥTs≜��܄�Rb��FR%�U���Urh{��@���L��Q=&ts�5k�8��ˉ?H�| W��7��yfR�%���O�,O,�]/*���	Ԍ>N�L�����6�,3Q�51��󻉟~t��{��#L�_|��/�ڐ�� %;�K����q���V �<����ToАc���Ƞ#�x��B���3���z��μ��F�%�/���X,4Ax�xԜG�ΗF���D���]��F�yC����
K�I=�#0�O��Y�>}UA?����@t;ƪ=U>&��Y�"�[%4��i1;�X݁��c�$�y5Be���3Q���T�1��L��	�:�)�"d���DsB����
s�'�5��U�i׿���I��'f��Af�y;�<y�L��j*�ْ�%\`�sV���m�WhH;m��öw���)8YO�n٣k������YX�S��P�؊�]�xwD���u�Q�۠FR�k�u	�Ϊz�fA�Lʴ���՞ꬋ�I�-�Af����m���3�� xm���G�|�	�<�0����db��ѵ���U��.]u�VvS
�Z�@X�INUA���ؙ�6#�a�ͿK&O2V3��FJ�a-��*دw(��C�9�Ț��̒��o8�z����R֊%�+$|i!,bb6ym�y���+��w%K��{�����x�[�>��$�ww�6�I�d���e�:�&���g���6,b������s/���Im�:mǔu�~2u��nDr�?'�@������c�\��VÎS��i�./k��L�0M�������A
�kt�<W���m�m�[���u�Dju�� �
�z�@`����SiM)�|�0�a��$9�k��z�H� oEu">������&E�M��Ă�&�Y>��S �'U��Fݎ�������P7V�8^��qT��=�A@�͂�zbo�_礪��lXM{�"��AFh��ۦ�q�x���w9�L���,1³T颴��X�/	h1��z�$�r�[�����+_���t��қ�OWx���K��������1��"�>���u]GK�1"(�x-�N� �h�I5����4?�e��l��YU�E�O-A�*s�1W�R���D�(6)�\�K�OZE� �\�O��I�姇l��I�է!E��؍�7��[v��:?��MkU��p�},�$:I��#����8�R/�(�k>35���!�	��!��& ����aK󝩃^��O��1�v�����[�#�
��_:gI��5P���$Sa��2ԖF�������k�h������OQ�8���m"�-+����sx�G�KŴ������Vx��?�t���J�Ѧ*I��Ns%A�������H�x�O����i�LԬ�#�_7�u�Xe��zH�G �XF:�v�[�,d�5�c��A��_W��2��]�W'O}٪$��f)�xߟ�%�t���:���T0KZ@x�*�>���/(|��Wz<�)o�M��H�3#�{�d��D)LL}77<��φ.�y���)�d��m�{�ɢ�A���.Sm�wZj�Tn���ic��`�鑎D���ד�ߥ_b_ ox��b�XlxVHYEB    fa00    10e0�&�
�|)ٍ�nk���ۙ�����{�~>�S�����du��mRM��	��:��EDT+շVk\SAF�{���hY;��KF�;T��jd4+��/H��n���k{��It5*�sw�jDD� �0(���>�iB-�{HČ�K��#z�����䋾�s�a��_��(U��w�'86�	05�t*h�6����)�l`-М���9��Ӆw�/��ۗ&n���f����w����3�	�����^������03(_Cx�~&�Q�OK�]�{Sq#���_S|�$����&z��pgv�ESУ��k�!���M�~��vw����S��C<��D���G����,�_���
��n���a�q�q�'����>��Y�ٵ����̌�_�)�'�����X��ȑ�LIR,��4Rw &��x�f��m���ð�~�_������q�������×�B��R!E�cx�xP��A���^%3�.�@j*T��������/�fK�����-J���\�L���U$�=����}.�|�uTEv#B���Z5a�S����+Ф���7����f���'e���Oa32DU���W�'k��^m��h��sQ�W����6�c�)$��=FL΋�N�j�w����G����!g��*U�� u��M9�碬-��1�8J!|?,��(�Bdت�e���nR~�'{9�����J����ÏU����X��a���#�����F� �
S�%��`��%7��q����y��}��w���;G�"�-M��P
��~�=�;��	����P�7.�[�U�j�B��Ћ>�nY���0|[��èI��2�vt���3���*V�:8���06z�\UD��yl��F���V�b_&r��e=.�ٜ2j�,����O����=z�*x����!)T�U'���$�:Ja�<�i(+�R+�!����_9 �ĐymJ[XF4�a����$'KGa8��Ql�/E��pxax)��Tǟ��p ��6�_F�5��g����)����_>Y����g����'5a/F�S�^���v�X��k�vV�_��
��m�JG�q��1=VF��J��ϗ����^"��U��2V�u{���˪�v��ʁ��W)�C_i��I2��)�`�����x��5dd�g�K�dH?}�晇~.�1ͼ��qϜڋ��-�Ju��e3��wW�ٮG�'<
��4�u�b�gz9N𙸏�Z�d�F�p��t%�W�� �zY�����癃���iE�V��@��0�R}[C
h;[��-a_6n����G��u�B�]/ΣY�s��5'���Z�37p��:� �rj���U��x3=��Q�aؤ7�|=(+LeN�%�s8�N�"�q��T_�a�~�z��Fe[X�ܚ���~����9�ױ�d�[p�#4h;U(qV�(y�s�h*@1�l�W�0�����Q��!0	}�ZB@��5��N7R\�F���x1�(Ҫ�D��]@u��܉�47i�Z@9����4*n6��Ab���%���V�14��7�|҂��R�Ŷ�j}?�����w-=�����d�9�1A�.�(m�z	6��Okk| ��<�O0W=�r����!�v<�=���ξF���k67�/��33Q�d�C�>�(2i�a�m��$>F|���[�ƙ�0R}UZ4]�
���7u@'���:��c5�W��T�+������XV}~���4�݅����U�U��6�v� [E��\�-
�:[yN����K�?��²a�� �`Bk7:���%�:�
VЫJ��#�D��x\�\�����d(*��4�;�,��]&Υ��J��F�ғ�9�P:��\?�~� �:��2.B农��,@���&-Xe=6e��!�܊*�f��:��ș͋X|�%A���\"��5%��>�M�#��i�}�R�{7�/�>��)�pV�>�>ŰCb��!k��g������I �G=n�Y58�O��c M��g@L�$"Y�1�27{��샒(����t�?})����?���'����:M�m���FN󽚗.��iA6�d0sOC���I�va�	 щ,<ď���82���r�SR���)��O�D�?�j_��q
�t�j.�#���	h7n�Nu��m�Ao���*Fy�Nr�&H���tpr��su�H�>'$���Y{��#�	�:S1��e��r�9(l��[P���~ٽ@��`VQr��<�����\֋�����B�ɜ0K/C�Թ�������Z�ĝG!B�VR�=�ƀ�E���M+�d@G��x87���un	�C�p������Sd�r8OH)�w������^�0��ҳG��UL�O�j]Pl'�k�T�d$�akY�C�$��K�h��Z)�Ŵ�+pmG�w�X[�ћX��zyں�=�֩l-o�M/֖�/�M�����w�y?-�2�[����#�S����oౙ^�7XDB�9P�S��VL������ � �%_8��� �����5����p�D)�������i��1�����M�='�DT8��w�G�2��7(��6e�n��[@�x�;�f잸6y;dH	���{]�@�=�e�����M���0e(�hK�f:���!Q+���p+(I��K����:Lr�(��+�:���*r	W������h��z�p�_������(S�Vh8�� �*�{�Y�+����"�VU0:!D|cxMvas�+�E��/�iTry��S=�2d�@��"��=�2�3���"�m�ͦ4\[��/����UR�h$1�z��S	3`u7/��� c���fa�����}8��?F�6�G�[�rb��ޚ�%�`f݉�Y,d�_QqJ���]�x�D���$�JiQ�`Ͳ>ߑIai�xP��wʔ����$DG�0!���y��C�
�4�"%��%�rꃲ�6�eݪ�!��L���M��c�+V�k�2.`���;"\I����^�q�8�mg'�N�\��̘Np���q����1'Cj�f�4�[p��_�s�f~�09CԴ�m7����U-�M��vx�vfl�O\dN�4Kk0���+���J���1 �t�6��W6}�D�  ���i�pw���Z\W�n	����P�.��ӄ�t��$h`�B(���C⦛�c������{�����&�<�Č�_�0d�� S4-���-pȬل�&v�ӯW�H��FjYj��0�����Ѥ�z���d��#����Oi;�?܂R1%�f��ګ��Jؿ_�D�j���nU�4�'�����5�Û/J�r?�����0vf��NSB ���e�C1�b�m�9,�c��iKR�(&)@��.K�Fh��Foc��V!�\��Rq�K�s��ٖ'����g){z�S�2>�wX�;�CDF��H20�b����f��������s�]��ekS�Ĳ�>�sL��u�cQr�&|��?׳e�䎦��(���:V�K�P��_�x�O^�*�!r��N7]}> �} ��Z���
Ӕ�3��IpH�ܐ� +�v͛۠審T� %n6yX��������iMUR�j��B�Yy��mir8e��o1]ʜI�}bA�
�zRh�uT���|�4r�R�cL�l���͕׺�~+W�P	�؆���,!:D�O�f��
\Ij6�O��PNS�-*�)V�!�+D�;�!P�t�h��1i�I`ҩ�����[��J�y�9
�Vz!�J�
Z�&2���ϩ� 
���Ptb�W�͝=17zU�&y7�0y�4
��㒿s����bgo�bC3��!�A�5�	��V�c۽��e��O�1�|��Fإ� �o����aű���S��Ή�:���R�I�*��V�\3�K���S[F�T87⦷b?n*&E-�(Y�-@�D���*�c��@����
� �� �D<ʳ�I��i�e�:+�X�8d�[���/�Ĝ>�� VD<�5��LPTX*ɚ�Eg*O^��?���b4Eu%z������� ϋZ����Io�5��w�O�vϻ��,�q�e��$N�?���&X��h�6
��A*�3�x ��G�R��!����K�PK��nUY`s/Q��!�X,�#3��p ni�wҮw�$���@��f��^���U[���I���P���U��%�ݜ���?��Ðy7�T~}���k�ρZ���o��4�,�~���e�D������m�L�������I�_nEP5&~�Y&�D��ݰ�^I$=� c�w�MXlxVHYEB    fa00    1860� r=�BܞPʧl��ŭl	Dq�'�򓅹��f>[��U�Z�Y��+�|�O`��!ڂ�h-5VM4�1\G��J�,�/��~`y�Nw�ː�b�x�i$G�w�.���h�4��r>��ӟm��h���
��nwq�Gw{d�U���	G��v��}t�2�,���2�n��1~W�Y��9��X�2��\I��W�=��%f�M.�{�2hD1����������B)'h&9�|C��G~�|Z�v����E4L�T�n��?*�°��6���\����OI��C	w��0�8
���G9{�	 ���Qn��L�����|o�w_�2��x�ǁ+��k�1CS�d�>⪗�N��V�\ Q�U4<������~� _��S2P���c*|�	��%������ƜqQ���^�g�S_d�,��"��TW
��J��O]��r�O��l�3e �]f���<2T��H	��w�1�iHD�k-���|3|}??�L;ء�G���y�
nc=���"k��8�)~K!�57�I�<�[�I������`h���g�
�Km�<�<^�.�@��sUZ,��èsԯ�;:��y���FtbB��WHT$M��6�8�Dr�����qW<��ιg?������������ӧ&��/�YY@/a��!��1��W��|��?��\X�4�<%���(��_�h;5W�ڐ^� Ⱦ�7�_��T����g8'g�Vt�>A�ҦJs�G��jդ�%�|[/�  ����_�E��F�P��ҫ1u0�4�"<�و���2^t�ړ�ݩ�ޝuN������7r[l��f���5���Y��RDnQ{�/����N��ɤ�s~b�z�Ti�sP�%�wnnD=mF&�ug�ƅUӭ�����~�T<f���N̏��??��%oὫJ�%o^'���`:�V=�)p/s.'cC����c�;ٳ��;��i��&����Ew�P�����$�E ��:��)됧���^b7��A�򞣬��	��
�2qo`�e�"���D� �.��D�*�R�o��9���K��Lg6���n�($�Pfkxz�,�v����gf�1�d)��'y��C������`/5Q#Z�v��9�[���JW75�Gɶ�K���4>Պ|��3$Ë��Y.Fl�t�@M2�rl�r�ˀ��$����_;�r��k��*�ή����d1����[�`ȵ! P�S(�Z��1hsr�>�'�ų?,2�]tO!�L�؛��T�Yb��E�Jp���-M5YT7ڈ4[	n�>�er�?�l�`���kU�b���_�e﹗���xQ%�-G(t��Ƿ��a!�6�ۼr↋�{�����*��L+0ZkĘM��"Z������e��s}��B����E"�N���mŋ��F]�F�z���������+�6B����O�&L�ԋ^/g�;�
�w�t4��Z�i���n�<Z���&Ż$�rpYt��2�iyE����%|ϒ��e	���&�j����t��6�j�����R)�|[[#�1s��#n_�b���MzP�7��W�_��*tg N�vX#�+�y�׀g.c`j#9��)G'0h>j��b�5�P퉠��K{ҩm;L�fZ�߯`b��BV�VQ�^;� J�M��a-�c�k�l,ޡ`��G�Dv7���E(�Q�Hȱ�X|p��oӬ���~"���8���F{�[�Oh����˒������/���ǩ��u��R��Ͱ��M��RI�yE ���͋hzI��V��SR�N��E4}�a�k�z5����yJ%n��������{��B�"��I�;5��B, Ǳ��y�ȹm.�ۋ�'�s�X�}�&[��N���[<��vI�'�J�	��.�Mx��A��!�Q�����|,F9Wȧ��������va�=Kt��(���>8EmF��#��o�y;���Z	[����>C*��-��\��t���4������k��]��^iȏc��HP�v�@"��[^W�z�G67��Uq�'z���y-�ŏT R���L��tA��И�Fӏ�����U���=OF��{K���	=�wO#�e��ߺ-5�F����r�ݣ�b��?rq���Wts�����8uXI8�铹�n,���( ���$�u��ϴ���:�������+���	��)�X�ݴv���>�1���R��%"a��ߺ��$��O�{��M��_�=��Ȓa]�
�q9x'�d�r���P6�xyl�8��O�u8�,��F�P�]k*�ĻPB*=�r���A�>�H��!���"��B8�`�fpX?n紗�d+��C*��˼V?��,��@�2+S�a�oS1�9EH�w �.��x���'d��h�/��|A1P��Z����Bw��/�+(���c�)�U*���Ft ߲1�Au�6Ms�B_I���*%�GN�j��+$�c��p�@˟��^�~�ʒ��6A��7dK�'I���ӷT�&*��9�}1h���l0L�8YWm��NG�` a�%6�V�
�'�U�a�����o�*�\�y(X:���X~On�:jK:�C�4���.�G?��D�V+{�:��
��	�O�16iR[���rxV�@��ب�щ{��5A�V�=-�����W� (���<b�^p��O�D��ͽ����������jI\i5$H�V^1�vP?��3[��9�'�@ȃ�I���/�_�<���L�Z:�8Ea�1d(�T����K���^z��ecQ�����&�M��@�lVۈo(8?cڻg�Sf�sMH��S�
p�B�?c���3N�'w��~���F�c����oBf�r��Б�s��E#�͋���D�M?(�8��V� Ր�)Jր�?}�GK�m�¿�;��2�E�/�Y��~�8���k� ����I�x������� �H=�<b�0�i�ʌԝ�6w{�G,#q��k'��%�^E�~bv������1	DRd�����߱
'<�+oN!��$��/g5�!fas��&c��,C�+\�z�SSjf�7 �Ui�~�����Vz�����(�m?�^(��H��p���ҋK���!dO���`w�w���p�ڠ'�8�3��mU������oFvD<��Q1����^�(�����bb3��j~j�0�p�M��؛��$W���z��%�6�[O9���`��h�jf,��p2���u#�D
ݫ���Ap���q����IØ�M��s�%�ß����!����g���k�S�ƹ�\�vp��^	��3Ϋ*B�M��(S.��ͧ7w�r������PC�oz?�,ͥ�E��}V�lb���P����ylI��W[���� �C��vh��YB�@c+r�s9evᖦ���|�����3%���[<��fj�/��<-r�UmM��J��B�'�(v��g��H>����e�-�s�a�#���{�*� "��j9o��#����%Ö��[Y��ș�03VQkg�G!���W&x�i#������IbԨ��)�;��n���K���L�f����`�a�6v�K�cD�AW 1�mUqr�*?����8U�>�z��lj��ߎ�KOY*�5��~�),6|���������D"V'���!�H-�v�U�qV��lГ(�=�ǜ �4��H�_<!C�m
����ட1|'���������J�����U�w��#��`~�
��.�����:�S0M]?�T���������E�F~�� ����z;�g_���k���f�N����|�3���4&0���3B�d��5��5]��zƩ��*/:VFҴ�{~Z�|�y�|��4��w�ޅݭ�A� )=�vB�pr�D�7�,���F�2EL0�b�Ȓ�� I`�*����ĳ��&,2�����*�\J$�f4�X��U�w/Ɂ�Bw�`mE��Bj��p�2s�k��%tH�r�Y�����X�e�D?�x"�Q�ڳ��M{=κ�@�@�U`����J#]h3��lbQ�&��
����X�d�9�{�Xb�K�O� �e<zt����t�,DW��S�É;Џ��:�i� �:��a�]4U%�h[��ӃkthI,|��"N��.~`�Ў�p�%�S����ń��M�w<�6��-�j����.J��� �l#�o��a��JG��j��?[�u3�ծ��T�x1��~eV��~Go��5A/k6�i�y������r%��2	�Ir�vQ ���&[F:eԕ��c~D�g��`�bS��a��~��#ꆙ�IZ�~(7�{�}���Y��B��ژ6����*W2�qП�\yu�0,�n�E�1�ᐦ���dO�[iH_0�,[j�³`��'mp]�-t7�>���%	L]ׁ���.?0Ń�����&?���~T��t�`'!���u��Y�B>��0خ\
Th`����zю�J������ӛI�;/�]��5'�]�$�8F��J�����23���ֺ�\�;�-�H�F]OCȟC�y}D?Z��J)x��;vT�s��v�s���)8��v�i �w�)��.�W>��ch�#ly�wh�P-�''e�iu:)�����V��r:7�6��9Sɨd~��k�c�=2��4���
�}:>�^��p����Wt~��'B�'�Rʬ��)L~+�_�~�Am�s|Ѭ�_	u�V��&1t��7���֙��������
��O�R�kT2�U���O��Y�'�1�(<5��g���d����U��k�T�y-U��y~
�����ڻF���"�����a�N8�3x$U^�-˅e�"�$��[Djpa�V^�K���|���>�=�p�Ґ����|�-���%�̨�i��)KV'��CQKQvql��?0����$��b(�ʩS�-��ͥ&�Cƒ���i�H�$h�E!�}0%�q���,4��e;�S0=l���<�����Y�C2��"���b���Wζ�����v���5)d#��	aA�Q�pK�z#V�m ��;�+n�\�c�y��M�6�W�2�8��֊FV��PN���=�K2BD����Y��d��L=��ů���O��c:����:c���d�:�L8S�G�F�FyB*+w�O2zMf��&z��|����0�a�9�z������j�'�2�DP��\e�W4Ų;hZ�ٓ���2�5�ړ�� /z|zx�n�5�dxzH�y�����fgs�d�i�qf����TT�M�e�\F�j<p���w��OQ����U��J���8R��\V���q!y8�~�:ݽ��?u0Pǖ����!�~��:Z���}��	�\����E0�HLV��;F�MןcPڅJ�%_�7��5q�0�a�8��A��dd�F� }�~̡F���ۃi�������2f����N+׀�_���+��g.�
��A����r�=Ny�0�' ��r��lh�T�P<�'0� ��j�;-d���M|Y����ELH1VI�iL=.��M��A#(��8����{�_���`^$�
�MF����r8�39(
�Ǔ�l���h!\�����Mv���	G���@���~������^��	�=i�h��i�q�fP!$��PK�-�6�H��"6�c��SE\��?U�����K7D>�g~�y���>Rì�(�*�/�~��	��n�����ig���	��G$�̏���uɢ'w�`�I�p��֘�q.����@�m�gk�Ԕ~`�Z�i�h���B����M�}J�}��7�n��@Vo��/x:�,W/R��B�SC��a��֎n���ˡ��~�BZ@��S�QPq�ӧ "A��/���I+��+��b�ּ�*)��b��2|��
3�MD=3��D	ɵ�d�ьQ�Q�� ��B��Q����gn��@'����oW���փ��
�uF�+갨�.J��n�AO�D�\|�2b�����!9`��}�z��I�ۧ6�@e���Q��P��6<��q3ik� $��р�����
;�bQ��r#/F��Dh��skr��/kÅ�Qh\���L��^�S�y��i}a��,;� V���5aR��Wn*�5�5�D*,8b��y��Ӱ��:l�T$�{�ɩj��^�՜��s��Z=� �M,�*�x|�{��3w[ڎ�-vVch,��HK���(�	�^Z�FCXlxVHYEB    fa00    1720�T9��ϔ��H��A�l�@�A��/�yUI�Z(�,���1nP�\VMg���U����Q�E^��@F/��!��. �p��:�:��< Hz6j�s��<�0X�
0g���U.�LbP��i�%��Ij��gT�T�ҏ(^�q��M|��⽪�mk\2�CA5���<�<�䃗nbQZS-�1�Z!?��8�)�����\�O�B���.o&� ������ZN5�[ҋ�[����K�V8���sn�����;A��ޖ��w;
Y	��ެ3�Xd�Z�Z�@d��7��V��؅��p�����x����fP�����<�/��B9*%}~�F!�5�ϲr:��Q��D���`��}�!ޞ�݁��+t�2<��׋��gRicB Rۭm��cQ�̻��x�'�<R���'G�M��<�㏓D�h�/2���d`^�j�4��g�	<��S54�w2��<�%��Q��x��y*;�=JMޥ�Λ��<r�_��ڏ�|�6�(���0��9qlR<޻t��Udz?K1����C[L���K>J4
/�>�����Yx���G'x<�����`�Ct���n�aE|>0{�H���ď�F��Y �K�q�����#&9�yq+��s�l]C��"Hč{ؠ&���)�!�c.��\0����YZ�%�����"�o��^�����XF���g��\{IPov�Yrtrb�X�P���/�)M1N�XC.�(�O�f����$���-O�U�OTg�� �}�w�M6��A������i��\�b)^��-��G�3r�4��m��\�������(5jR�hU9B����G�6(� ,[{���KjF4߳�8������Eьw.|k����&���s��e�^i�'$pS͓%�)�!ݺ}����jGO͋�I�89��a�w�W��{H��;�kX����r�{�X��=�h��C�Or�����b����AԈM'�#����`k6f��8���� ���C%l�L'�$�|q�Q�M@��}_�͏_�Ҿ|��yu#Iu�㣂��@w���j����D���E�.��h��ra>(���)���̋r=��ˊ5���z?��8ԡ��ٶ��Ϟ�rn�֎L!:&_ػ�9G9��+Ukz��9L���c�ӱ��{yJ�9�^�:1�:IQf�8Z}���RK�q"c�z��h���V�7B�����r��l�K��h�vՕ4�<<���t* �ɴ]-N��f��+��������3�E��]M?rJW�`b�S�E�8ze�����.���R1�v��:U(@��ݪKJ�޺�����M���]N��z~'莎!6��IJ���BU���M9#����3�C9!��DXt�E`�b.���犊n��(�9����{�9D}�4A���U�������3�'&`;�)���)'�mc���i��x��!'O�[��8@î�zUPeW;0��3r8�$�IF3���~�l;9@N�:�����2q-�w�^b�����O� 
�^f��'�x�%��+�(eMTt�=}i�&=^��;[Q=$L(ae��؅5^��T�Tׄ�V��~�#��z�_�H�E���=`�!�0d�G���~���mYt y���D����SP"��z��?%,g@�yB����� H�`f헋`�_�5��w�R>����/����%K��d�M���
U4�PH̫��U�'�kQ�����2G�/��4�x���]oq|�
E���3
�#iE"~����U�d��:{���D�JX��X�R��������"a�/tM�P��.�� )Bp�sN`h\J=��5�ݬ �o�_��	g��Ń�yY�OyZ�)"�*��Q�W�����4�6wg�G�����涴�Q�m�V0��Y>�0�?�q�Q�	��q3G�p��j(ٍj�~$���7�I?zY����Ny�C�]�3��t~�긳��֋����q�'�2����?d6қ�7NX�]�A}���^�SO��Q�D&�'�L0|0��K�o���q�� ��2�A��X4��f�ш�������6�e�-棾X\�8S�<޽�{GM����5�|�<� W5;������`-�%�N�N�!a^1\@|c���r�z��8;��*$�fR�@!b����1��@��/�m`pi|�n�n���L޻*F��>s�O���ėJ�����H!��/��ޙ�?݀�C��o�e����أѩ�������Ĥ�o�o<:�r��p�9#����[^�A���&��o�/Lc���.g��7���2P�Xx�ƽ��Rh�R�%�����;�&���� ��Pn�$�����J�]el��=@�h c/�1�ES�o<V�]��H�������v&���!g�t���q����ޕ퍙�ʙ3:D>�D*!'y*��j�����䣣�ZyU}} iY�]UQ��X�ҁŭ���7s]S3)*�y�/~]:�Љ"�4��l��.CM���gS#�̜x�Aoj�	AL�������(^3?���j�B��! ފ����e|�bJ��0�����c�X�X#O�M>`���TWaCՏ�_���V���AS�[�R����I�C�I�	����t�ߝ�H���a� "-.AX[����'�Z��^r�dR�e�$�U�,%�u����8���YD2tz�/ɳGZD,�ħ���l���2�7�?p���Bf����e���t���8d��k�[�nGnoI��S	�0W�]'�/��]�U��|�����[!�`l�Y�F��yr�
�"�4�E����\�"��뚿#�u����a��Lt�6��8�o�K�K���<6�~�^�j����]Y�9��C��ϐbB�L��I���d�o����-�#Y�}����P�-�����S<b�u�|��$Þq1��#^��b�c�F�g�D������m���d��^������u|�y����s�p�1���&H��L��N���<L�3 {���X��;���x��@a�0?�',�h�{
P�	�����2�e#��8����Cq�Q��x���_VH�~���Ƅ��I�(nw@�Vq
���+"Z����3�������*灻�P��Е��O�����^�ve~w7��2Ig+�B'�Y�I)�bb�$�0�=&��$�:���{��	���/Xs�xg���^Y-�|�r��i����d�k�E9��4�{�?�씅c�
���h���|F
��3�0�tq�~[�8f&ŨY�ͫ�}�7S�s��e�0p��}�hg��̫�K�d�=���R��s�т�����h�v�=u��A?�a���������2���m�&��ĵ�A�V�sV�*t9�C>�D���S�Sz�[ѹ�^���!OO�
���?Ơl��!b�܉n<0�W�drmOD+�>���b��,�T�~\�g��K0><�ҨԽj����v;C!��qb�ѵN��z�2�=*�Ո�]�����8/�`����H.vp����LJ{�7�+>%DL�D�C)&#n� ���2��(�-$��:H��z�"l'�'w�g�?��w^�����[����O"29�B��E?>`��t�����~ -��xI�Y����Y�%�:���t���n��ۍ=���/�N�b�6�h���kZ`L��A��|&R���(�b���x&7%������V��	9�'�j�1��������`P��?��]�	Q�A�A�ه�gud�l���b�LT�����5%�d"�����A���v���cRh����@\�f�M���D+s�^T�or;�1?r�{�(=fy�_�B�N6܍v�Ee�+���h�2�V����U�谹�,L�+�O�i!�g�	�k˺TP���*wZ��":s��»7moe<��{]9F��������T7<Q -ö�UI�����5�&L��C�<�A�EH�������ёw˗�����9� �����q,
dOt,��ا8� S�~<Hɷo�3� �W��H����sU��.c�O}KSfp��(���c�|��˪�E���~��<�=��Zÿ/�6ܬ�:����=��HLZ��\���7�V@Ѭ�����m��n0��/!����U~<H*se������{�p@^�E9==1���^�����}��Y崛z�ټHͩ>���
�P?�|�� l`�wS�MQV����ٴ}���f�;ر� �"� �������{��� 9m��(D�}9�C%.���V[5�901�§f��!��@�Bd���;�tG�t�ϣ�H9�P�q�˞^����&~~���	�p�y���J�G�wj!�H�<J��ţ���g�����g�U	� �5�����Z���8�.8���3��(NS�������Յ=O��G�aa�fi<:"���Fp�
�Wbo�����;>Xb&���v	'?�P�_����T�S�L{���o?eS�(��2)m��Tf+�m�҃���>���`)�)w���Q��2U��JͿ����N��*0ڷ��KM8�O3b��MeKj��W&;�٭q�?}8z��T��'K��`����,0��L����{�.,���6.\'��;8��L
�@2���3��������3�o�T�q[�dY�ɒl��|������C2��.��6T����$�=5�������LUni��?K�M8%�\�^��>�]�H�]�f�cv<�� 0���A'uR#��It{�����IC��4��.�����1����a	�Z�q%�ѻk���5�2_�Y�����3Y�<�OI��}��kʞȁ6VN��ք,l4D���f9󖘴+�'�e� A�s�YkT��gI�<R����w�KE���)3A���V����~�e�����R�VH��FE���d]~+W��z()���fQ��G���v����wW;)^��v��Nw�:����_ac"�j���B�4j�@�s`G��`e��?ϲ!5�`��s�	Ep@���Mhnu���8'���I:�I �����p�����يh���<��1N�^�ii�N}���N��8NQ2�桠��4�.��&Z����_m�~������p��/<r��,g�Z�	uZ/ع�T��K�<c�
��,����%�&ܟ����Vd��њ�k����?�8���VH�"nY1����� ��2�wo�H6c�?�����n���Wz��i��IS�
�7ۙ�$��l4p豋U!	1���~�yY~�E.^P~���^�W=����E�5\��+E����<�Jӏ��V�����`�E�J��������پS;9�+d}�g�$J�^y�&)Z��<�����4����}H��zb���W����MY���"%ʭ��(A�LhH�5��s$W#�1�Ɏ����|,]�b�o�����}��6��h���(��C��T���~�<��m�C�Rt���8�}�5��R���ާ=�yh���u��y�HV ^���Q$K2bp��="J̬�VxU!�o��\�;�b��BJ�ɍ�#���m��%���ޜ�U�L\�r��a�bS�n'd�Hb^�@VZf	��}��sT�~\C�yO��9{�� 9�*Uu4F,�Om�OIio��d��خq4߃����Q^�,���l���I�9��GFk�x�_-�����~��bs1�S�KEDk>����YF���$�v�Q}���~��ӌ��u���
e���0��F��G[��_�+ 9!��V��b������0�]������Ck��k4=%g�*�ot[z���1�������d�rl��-�x�Å"\m 1ϫ|�ŲR�蛝�Q=��v%0|�}��E���7�r��ҧ­XlxVHYEB    fa00    1500�K�ӻ�J-�·��5���6�C���&V��j]�yŧ��0n:�8&��8'*,Ψ����/�c��
�s�ؙȚ;~YgykA�sUg�j�C�Nx����~%o�Mପ����lz/�nz]���C�nZu��y"�F#q�K���b䒯�)ǯ��м&�S�J�J��ǥR��om��4�ֳ�M!h ��;��q��r�''��[x��`iIyQN�x&��!� ����El��3����1���D��?�n��sn���+||
]gx%�Z��j��1Mʲ�/��/`���m`�����d���q�¦��EL�#� {�]	T�Y�}��q�z�����
�l�Q��X�����p'Bl���2�җ[�6�U	=���kp �յ5i���ON(r�|���6�N�J;ӝk`���W�����qԩY���\�)�4�JK�y'y�	����4�C���;m�Y�E�o4�#��r+[ь;��f_���`:�h+e�
��FO��^L�;0�In��ݍ�u�ӕ�e��QZ��c�����p��X#u�3�$y���w0Ĕ�ΥV�'𬋟���Zs�P��j��QZ��S"%s�d��!H�V�k��i$-��p�ԝ���N%����6�$7�;��nЪ������r �
���9�$���DF��^��,��3.}�0��[�!�Tz��ח���N�5��AI5p�rSX[�񢲵ETҋ���#9.��#|q>��D��O���~p�C�~��;#2�	M�5y'qݥV����y�+}�T�V�ӟ��+u�;��Gf�"! ���_����j�7(�eFx��޶��A��4��4^����9eW���5y�L�/Drb+|hG$���1ݙ��%�M�x�5�J�8��f���Y�����g�NU|��Wc��(k�]uء6��4lX!�4(lZܑy�= J�V�Dʵ�,Y����c\�%*X)�Њ$������ՠe:�'1t��T7��-Mx�>���4֓m?���Y/%��4ҝ1%`d�����dv��e��rI�Q		l�L4��_�9s@����{���-�TKnI}�er���Tt5��M��i�5e�N�Z�+s�pಂ#�ƴ-V�
س���O�LQ/:�'5:��d���i��$��v���^���|j��)� �B
�vX�}��q��y*��st��J.m�x�E���U�:$n��k�ո�;��¹<t �Ts-X�C���pT0�j��CLZ�'��p.�*���V�uH�^߁���6��H��~�F�|��Os��JT�BV�u������J=�ޠNF�d�+�2vP/Ek㺄L�:�bՁ���Ȍ���ve"Xl�l��V&��rD����u���1z_�aL�����j�!��4��������&��EQ�G��S���畅�o�DR�CU�s>�Ka�=��Z��@�Š��Y��O=�P'�ұb09�]��;��� ��|SvWY�s�Z�!��7+�ګ?�-	0���(�c�Q
W;o��FQ��J	�R�JJ2b[���*��gA[�\�b�� �_<�kF�*����W�-�;)��U+�:�U8o��`&�(���.���� ��Z�,۴d�D�J���m�^���dZE���OnJqϓɶ?����Cy�P�=.^lN�>!�%���2V��'�9�~��o��c��u��C�\�J��� 2����_S�,��h-%�Y-�ҧ�Z����R׸���?)\`�M�&�Y�y59�3���O�<+E�P�z.�$3/����"N�?��F�������s��k���u^�����:�i���&�<Ҍ�VYZLP�İ��G��3�, ��Bĥ���ۃ�o%�D�(�W��&A�_:?��$j����أ<l��n.���f8k����@���#|�o��i8POy���!�N���<&|�_���ڐ-�9FW�
!�%B��腝pٮ��#�9��XNy�Nï�Ǎ���/#�G�ػ�E�gkO�\��)���8^ڐ���i���4\��m=Y,��Fu�_�|-�#����j�R��o~��z�Pi�ZX��W�>�!L��0'�L�����qե�P,6�7���7%["�8ٕG] ���S�m�������Y/}��lZ�~�c|���{F�J�Ld�cﲸtUӑ0�ma�D�K�D.��s8���{�rh�Q��U���������?�:��h�G��0�����@�����P7�ݾ{���2�[���x�3���Ui݂���5X�F��Eʈ�{+��ߐT^mVڪ~0e�Wz �1C�O���U�U��\C�r����M�=TV����j4=����䈫��G?����)-�魦�x�k��o��]x�pn�B�t�H��	�|�8���E|8�%�O)l�Ǹp��E��K=�೺Z��l���r#�c'����H����/���w1Yh�Y_Fj�?pę�xg:&�����a���f豴����5�1m3Kl����u�D-GR�B�i+.��	���;Ə���������xp�]+�Z���zDв�u��{�HY��e���oI���b����CVZ�c͞��'��#j|�P"n����f�&�J|��v̹�7Z��~OՌ�~/�7���.k>S�})-�sJLT���PRBkU��K{.�ED���?�k� >m�r��I5j�i{إ�X��9jV�0!��5v.l-J
�T2I�N���	����_1aqw0!K��~^��F���s��s�|�Q�+��?K����T�t�����s�%]�q��)*�u���٣�I�R�����:��C�3�j�PzX9+��[�/�*Z8�
����+�%8�ժ��γxR.7n��E������6�� �Ƿ!g�	>�b�8��v��^��@J�����-7+���j���:fE���ɬ/U�d��T�7������w9h�*�>ʌ1��PT�����_���cYD�ڹ&O�j�\8zoM�$�Q�$qw�CBwՂ-bǇ���h�]}p&��B4j��= =������g$����w"�]M�eN��}JF���Y#�z�dl�]ăɇy�â��
�Z:�g��Ӎ]��-����Ȍ�s��Μ��d���2��~�L̻��8�����46�v'U�'8�)p���0��/��	�㭉P�h��Zt"_O�6��Ր6�a"��S����'f�h�-Df�(+�HJ>Z�ퟹ�x���~�}!iS���2�S�$5`6R9��-P*}��+
b�6*2�WQ����J���!�h�l>����JW�8
�P�B�����aY���tm>�T���
�B�O�������Sh�i�:i�YUk�γ8s�D@:�|�ۯ�t�~9�M.���`���*��8?w;T&��c�28�^C�D�?X��B5��ɇ��a�O�iΎ�1q���_l.�{���a�ȇw�,�� E��`%�y��Rև�ƿS��o=��b�#�T����Ka�질�����\����1�Hi���>�&B鹣����Gc.�Pd���O�`JP�qpM5fj��Qݮ~.J�����Gڄ�]ǋ��:It��>_S���Zj���[II��F�%�IģW�� '��:Yޝp�, �6�|?`" j����﵉FՄ�Q�p�B�S _տ	M��9L�"	D�ꒇ&sFF*��	�t�њ�[?���&�&C�]˔7I��k�{B�7��]��%^oz~`AH�sr��c��+&�浇�
i\5�;�/��,:�^;纽�&��EW�Lm-��o�d��ـ�����f�q>��"�e��(���nx:�3�"�Zu������?W�7׳�W[���z�Y�Gb���*u����i�Q-M��k��b�/p?�a���+TY��?	L9:֫I�倀��&��V[V'2���[�@���%3�լ���l��{)H��w�n�����W�=aG���+�w��n`29��@�=R�0��m����f0> X�$��f�ØQ��1`�JV��2`�8:�����	K9���H������%�"*��iT?L��N'ޖWlO\оBt���7a���꘠6$����}oO���3��x�F��qC����E��G��ܥ��o�qb��-�Jщg���~*fA$CGV���헔�y_M7{
��d�~�� ���@�w�]���7m��,�'p^�Ywaۋ��\�x�͙�Z;���Y�=�Y:K���g�3�Y� 3P�X`O�&Cb�C�1������W��|��ZD�ʶ��8Ma�k=�n/�A� �iZ��D���D��e��	�1ϧ5�E���]!�F�/��p/ď.��I������K<�m%.����ձ$�ܓ�y�m��:o��뺦�p�R��k/���C�.�O_������JX���:R����4� 1��#����`� 
��$������i�U
�bI��&*�3���ƈ��˯����U��ђ�{0[���Y�W��Ǹ�ǫ��/��S�LUi5�{rx'�b�zA�J��M��t�G�[�c�PpyF;ܗ֭��ʁ�1�7�=/�H��6�N�w�X�y���Í�|_�#q�YTi��k��`2���2X�n�����(��K��Q�>%O)��Vu;�$�����uwI�n�'s<��5#�a0�繦���}Ĕ�y��T��BYW�X2 D磹F��8�B��ܱc><�(h��������q�}�kg�YFIdmg��m���"�0;U!d�ߋ8�p8���6c�	-#��N�Д�_o���#E{SIh9���I'�no
��ȸ��[�{;�����Aq����{���'ސ��{�]m���WPQζ��<�uP��s��V�3pn��ƻ�*X�H��N�G"�q��lv�'J`'�<y������-�L��������{�m�ey�L
���˭lG"�Gr��\��{YE�>�p=O4�#����1)В���Lf� Ұ��W%�3\�{j�t>�r�{��HX�U��%K'k���I���&�މ�3*�E.OK�3���l���I���j�x�B>Ձ�"���ZwJ�wc�-g͟���j1�+&����d�}1�䬽�Ժ ���D�x���Nؤ6��4|�Oy�ԓ4yV�*�:K[}�/"x�����v�}j����Q���#��#�J�,�;�+�Ϡ�hLΒB�$nq��� c>��{ cXF�$`�ᴱ�6x32��x�(��	�p^��s�mP�_�|<�Q-���	:oP��arb�eeS�(4f���)�Z�$J��7t����0����k2��`��t���XlxVHYEB    fa00    16c0K�U��b�|�/vl& �'�"�;�c7���fs��rݠ>O�b[\!�HuC�����X V�ol�mM�^�H�~L����)������NhX������[�TY��h|�髸��O�����K��Pf�?P�`keK-M�g�و�����]�W"7�̿S��4�JU�&�:�+��te��Ź�7���3o��D��	��D6ϙ�E�h����֒��#;'�� ��?�����+���J��ӽ����ƒ�ցJI0ژ+	��TiB8��oK��ψ��}�k�뀻 ��`{x"�޳�b|��%��WL�-�1H�A�hk\��^�a�d���;������Hpة���_X�����4��}��#�ȫ���C	̺r���ޡ`w��KS�r�mD�n'�R��J��y�WVvS����%5��㩟�3�� �q��-���i3�M݊�+��D��SaT��L[��C����Ip^�\�<�L�{MD�
{Y���\�\���]�a�;���j �x�h��yժMjR|���w�^��CR�W_$�t�!f�G;.P�-Hc>�.��kk�>��>�'.I�0.��6jh"��1l����\������L{ �:w=Uq�����٩߶5)����^�M<_#��*�y��@�Q`�?~Rk�[�?�������E��?V�u�Q��ss����hꛊ1z���J�l5���d�\?ݨn�_c�N�y�[�x��r|jK�5aC�Q�/mD��(��nəf3�\p�j��MQ��٭�ДfM�����y ڼd����udk�tha�9G3< ��yݚ�>�-#�" t������������N��%Qx_��*
~oրMw��)�d?�/E�»
�_���K�U�f�(+��%ʾ�}j!H/���Q����+�f#ډ�k xdx��Y)%��{��~���KS����+��ѻ~5���]���Bb����t��ڣ��^"x��e��p�R��\��I�~B%�(4j�G����(!*g���0!"�p~�gmX�s�e���vOB��7���#�ŭ{ӧ�o��O*<I,�)�<4��yn��k�	4�U�����BL�Ӿ˶��]V����N�(ʡ��?a��׻2���
��v��2Y)�|S�*1-�L ��Z�c
�JPlz#)&P�������Ž�;â��H������M�{CA7>��llE�^9���X�+l.oI!R)��?�����z��X�_CV`-�N�2I%heAz�gB� ��	��{����I�b�W]�t�����7�\T-z�v��t�� ո��v[��zw�fk��Pj�3Ե-j������z����+Zk�`�:�<�:�� ��h}
+*���Y�g.�z�9��H,mX&m�Aա&Kj����{�&�D�2>�|���X=?�M���KMo��&'t[�����X�I�y8�:b�����4J��#A̐���R|�ˊ�faB�GId^��Bm�Y�loC��Z���>4;Mz�Mza���
�$�f�J�ǈmS?Cy�e��Ç��\D�>YGL�~^��Jm�8�X�vhZ�4���H�m��@��0)mFd���U-q̣Ҧ������������h8�x�1�����T69kf�H�QA��B�DEyDc��KG����[$e_/Z�!�����KI0&a���r�>�(Y�P��@��a�k6n!����؝+�ȻJ�*[�SLfz4��E�������H~��(sbT�Wy�bތ�3a�.����L�\0�N[�3J�ڻJ��e�̓\�����_���)�@�?�Q�`�^�Y�1}��7L�O$NG!8"1��˸��'R�;���k�� v��ψ�i؍����JF;nO�k硷�gÜ���8f�V�%��,�	��\�fʓm<��#l&���M|"�M����G�	�Ns�u������C̅`h5�F:C�:u�O�m��W���fpPP��bM���o��)����V������w�M��Ԏ�AA�ĭk	����9�'o���J�Bh���D�%�O"��٥��f�]�ץ�Iߐ%<w�F�i��o���w"W)�	�~O����i-��v�E�b���A}�?^��Ř��ܮ1�����o���J�m�]A�fIt�}��X�q�����_^�n�t3t����7M!�{itL�T�Oq~�����w�D'� ���h1�i���JHr�
��qy?xݽ2�2�ӄ�6k��ԊV��r�8��Ts
���|�۱ƞ|����)��>P�.O��~�A�"D��ry�p6�16e��s�Y�djCS!I������c�B��U��l�t�S^Tq�%A8�H���[���[�k�_��:;wF>x��d���;��6ܟU��u�'�Ť����W��P�i�d��� 0r�hG���PVT�H�E�{8U�y/�h!��9W`@;!�~�h{���h�P��.�j�t씏mH���@���tk�#
�L�����P��Hѫ}�4�4�ݷ5�L3'��?3��g����wEW�݃��h��R�Z���4"P���:;&�7eI��d?��Ќ�BT ��7c���X�z��1��� ؇����wuܽ諽��Zx>��C8h����(��SO{��׃W�%Q����AY�-J�`<�����n��/�D�%�HWI�,g(��芗�:�a*T�h�3� Mn)C���%�#}ߧ�n"�S��0��r��E9L9�RM?0���=`�$��M7�@�ZidCϸl�o/��U��Q�����E�9L,rr\�D���]��Ƚ�i;�`����X姺q���p��^��*{�������U-��~T;}��Ǒ��@; �a��?_��0!��z	aP��X�e/y��e~#�G���]H�n��W ��<��A�	���F��~�~Ҷ�u���7�gT9�j�7��݂mi�JƠP٘1�K��ՅЄ�]�?�a�-���{W%����ӗ�Nc�:7�A���,xV��ALPmRg�V]Kw��3+k+���nȠW#������}�[�?�E6x�N�L�|�ؠ,�Ԡ��UiZ��`�=R�i�u�M;E9���1J��
wf��V��w��P�I0:TZ��?�F�[�7e�:ia���F�Ho�X�p}߽��O�	��a:���;w�(��#R017v�i^�D�
U���2�;w\�%�zD�_�N�5��N��HO���*��덽����/��^��h�I���U�GYP�*>��3bh��{w��=���-M)�=�r���܀�𨲉k{��r=��;�x��gP�w��:��ު��:��6x��
�Ύ�|@�y�V���Y��A*�_��0�L�5*$�ۯ��)g=�P�*�m���!��"���F��f���%T���e+Dz|��1:KD��B�����h+5{%�:M�S��Vf�Gd�55r8��F�q7�(}֋SG���
KҒ���9�x1cp�69���S��q;�ԘwiCZ*ZQT1� |u����Do�� W1;,�Xr��zz��$���9�/k �4��_9B/%��<M���z���9`r��}v�D]���<�~�q�)�(�ۅ۫�
���o�4������#\	�|�
�(Ő�8kb
�e���`��SK���h.Q	��k��Kj��K�Izn1�0:�z�zW��c�H�l�dc�adeO�\�8T_N�P&�kY��iV�"ҩ���ձ䈧��i\��簰������OWs]l���xo�bv�-F�\^F e�8�UF��A�b!;� �.����c�Wه��0���r�΀B�)�^�,�!w�9 ���H#�忮��������[\��ֻ:�*�Si�a����+�5�ہ���h ��_L�c�7l�8��Q��A6߱ ��'�M�+�[VvcmW.:D� �%&]�ֲ֮p�����&C=�(�Έ�^=�{5�
��@P�e�VV���Aۆ�����$8�e����q=��E�5=����WŷFs:�U|�����'�_%�F[��Ǵ����k��͓�M.ItZ?�&I����wJ�o�1�)}�67V��=6�2+7FH��f���ԬÝ��o���"�y%��s�C�]�l8f���t�{���v#MXuU�h!q�'Oފ��S�X�C���F� ̉��ĬM�fHf|�C��1���3�@2g����g��)tH��	�,L$  ze���!�`�"tO;·��\�)8�|mf�����u� ̭�o��M��mv��l��2]8����3тZ���gp�N�)w!�f4R��)m;��0�ˈ`�G���׮�faǗsK�@~�=�v�+@DAH<���/:�TFI��ͣĺ`"2�?#�XT2H��t>�qB�l.D;)C�B������cF�ֽ�]iW,�,T�z��������)����:�����:�,Q<SOw]�2��v��?�#���o=��8vi�W,�`/u���L�5�\���/�y���Vؗq(�%\� ���q�LC�.�
5��:�>≏5f"����G�y��v3C����x��e�[�����h�٩o��?�i)�Ě
�q���$�	yW�*q�3������������j��`�=E��v����%�P���\�I������^kq1u�M���	���v�?��5�Y⠛� Zb[�n���ꍟa<�?cn�ṾKiU7E� nH?���<z��U4�7��{4q�؛U�^+�W��a����ɐs4l�ǀA��] +�x���|��儡�%�
�Jv|��E��Ta���!�� �z�J�=��Fȿ�=H�m6`�6H!���^��Z�%.\8n)����.�cn��K_��x��>Z=��~�ڻ��Ψf�P�� �  QgS-L���x0}�#5y۴��qiY�U�[8�N����M�`V�-h��ޏM����1�-%�Ѷ:A���`�sk���wC��%�������$��������?��A���*�U�G��J
_�_��o��7u�{�Wc�T���I�1�a �*�X �X��i=
K���9�p�EV����J��^�FJj�D���#d�ޱ�"����q�*<����_���A>��G�`�;5_x��ϲ%ܨv�\Q�Jy��P���T�d�f_H�0�S��Z��G�ͅ7GRo�v=;�����B��	��[�S�p�Y�ý�j;/r���pc_{��0�sp�J>[�������F���]���n5V�CJqY�yb�0\��X<�;�W���0د­�(d������(v.�����H�z�.���ր�},�"%Ƀ|L	�v&'�2����kDV�>�
�'�����@Sw>�Z��,�E���u�Rbii�8zFД����.X��Ffs�r/K�Ι�8F�P,ns40�)E-Z�ܝ �H,��-��=J䞾=I���/Mw�Tѻ�6 ���y�vH�����
0��19a|iZ*��6u8�!_��B �#�:�JOR���cW� �(���W�S��l;�`	q{��ۂN������2T`����������B���,JHic��]�r��y�9Mۘcd��з��*M��%�k=����IXK��S��"�qi|	�p�'1���q%��D���WgQf&h�z)|1���u���m�Z|�Vg`X��6
H(D��l�(s�F��w����F@�����}b0�\�sˮ�mķ�ƌ���+E�n���5MHE�JxhZn�7󊙌P�wW١�B��Z����'��zXlxVHYEB    fa00    1740�i�i:XoJFl��� Vq_�b��G��H��d�5�ri�昋'�@����O�B���1|*?�}'X��:E��BXiۋ�c�������^')x�h�y��Ѻ���|�1_Q�6��ϋ��B�P�^ȍ�=h|~Us�gS��#7(p�����IN��eJۦ�6��ۨrnП�?R#B�s!��	��La�5��3Tl�(��W']|�2�������)�@u���Q;�)��A�xuS��K��@����F��^>��(,D=8���TxC[w����;r��H,��PR�9���A���k����en�A:� Z (�?y5��X� wLQO���ώ�S�ۜ�UoNe�dݖ?�� M#� M9+ -�[1�x9�O�^��?��"�cX�U�FoIWK�܄���bm��$�b��(���9��'�C�[���+r��eY�nf�*#�q���P�����= �h�B�֍��3j,��!Kd��O��D��M��j�\���g�R�F k�ג��Q�L�8���(�֘ܜ��Õ����n����2�u*
k�r�xej�>C[����B���l�c;G5F��1����x���j"�d~R��k��������ҳ��T h�}�x����j�<q��-(����,���WK����f���%�����a[�#�Y
���HfJ|j��b6��Q�-�έI�1���QY�K�x�8d
�+o�Ay���1Y��e��� �7��[֢��R����n��z�v?":U���|�%�aS��U)�����ދM-o���TH�aXu�x*݉I�����L������
�-<KR	��?�<T�X����룸�S[Z���a�0�$`���q���Nɼ�B�j�#�"����h�s+i�=����Y��.�j���Sбv~(���#&9G|�)���Vϱ7���7rv�ǵ Ӗ����
h�A�Y���u��e����F�'\�֟[�6߅��}q�*)�{�������k�.MQC@Y�#�wW�l��oU,��؟����jEO�G�!W��E��˒�F�0�f�;���y$M�j�n�M��Ō�>���hF�i�M����� �'��xN��9�B\@�����J� \q�^���0��#��J�]0]�,����cy��ԅS*�3��1��X����m��K�̽[�A#�G�>٦"�������mK?�A>p�a���9>��|4�� l5s\�OJ`��"@01��/�ܭ���j�{���ZK�*-�\8��z�ʟ� 1ue�Ӧ�JϬl���hq�9u�ćUh��+(��>��,�����������D�pz����U���&V�z������2�p�(K����i�������g:��fvWj9	�?�|�_qx,OT�>��y�h�˳,E7�[+�Qm�"��=�8ش��� �;��I{jދ�?Jf�Mlh�T&7*�+�L���U ���7Fb�<B�GEP�� ߑ�DnKx��SrƆ���C�3�$#1�l�
K١�z�'�AbYȳ� " _2�����	�j:�kD�Cn��z�:����������8q{��Z��O�?���f��E���1���@�'s٘���`T&�]�JH����j3�)Z�m�����Uj�����̿��,(��"H���(.
NQ��dc�A/���;��G%/ ڳ�%�=���}�0U����4�� ��[�|��\�"��' �֑@�깶������ !�}tNo������(��O�ژԤ��C�$��Z߁����\#��Z���/��[g'�@�תŊH4^���i@��"?/�����c�t�z���/�R4J�Aĥ(_����)紇�]$�a�t/�HWl��B����a�n4 A�
��$�n=9��H_��!��V ��R�Jq�A��q�,q�I�������f���=%}j�Z����As����}Es�Zw&:����$�XI�aR��	3�v�M��s��G]פ�`�RY:d�@��a�#ߍ*a����:�~���I&�jޓy�;s�ҫ����S)V��L��G���BM���p���<ȁ�|�ڷE���j���z#}v�x/ʛd7j1�O�K~�vh-Sh!��=7&9�,'�]��f]7�tP0��̈��\!3'b�~��?s$�Y�հBw�i��<`����>Tє�%#�'͟�����C�?�}k����^[N+�(��b�gn�p*D3d�gP���i�z��|t���J��z���0���c���@���<��ť�Rt>���
��ë�S���7�ĺ8�ϙ�%'���~5Gٵ?��3?%ILb�[��R��k]�����.��(5�a��{��ִ�����i�c�"2f���{p*Md��;9�F7yQ�hM4�k�)L���Gg6 ��JO􈌝��(|�3�	�Z.�fN��^�۴�DJ+e,��~?�؀N�o�{,�/X�3֡��ma�4��r<fo�J1�{D�>Q^�(�J�2�:Ibs��Q˄#!�UB��#� �%�|���ʦ���\��M���J�&�楾�B{fD�8�2 ��vyx�t���S���`#�'��n��UB�C�T$f�~4Y-gek����cuu.?d��\�xf�U�DK���B���gl��̧�R��θ�<�e������¾�n-��s;Ү�4��S@UZ�v3;�_��h���
w0�mM�נ��Kw{��̗N�I(���E���ސ�K{����]�*Ec5�������;	@?��4��%�ȴ��т���
�:z`7�{�b���@OaO�IzM(%��Op��Jc�M`U7t�����WJ8kB�� �}���n��g�׬:#,V��9��][L�H�Ml����ؐ�M���N�f�V��^v~cu-	��&ߜ�E��c��J�]��P�g�Ѣa�9��׼�OG�1,��r%J����#A;����`�z��1W�-ݱ�����x~e�͝��3�tN��Iu.�W�֔N�|�˳���)���m�|(c-�E��P����B���)��Gi��k�=4�6��怗�+lh���1HL$�H���+��,K$ks�ŕuv���E��q��r��<��{���a7�+��ye��^�WЫ&����Vu�2�ʽ��ӳ���K��{��@I��������8̠�
��^c�]�Q���B5�bpхz#��N�I���⒚l�C#�EM�>��ƚ;�(�#uU*O���E #��@旣���E��9��ᑮ�E:FV��m�BG��X�W����	���U���[;;6�$���R�4�rP�w�p�wo���� 0<��D �.����8���Ah�,�9��t}9����H8��a�b2��,Ұ�| �ur.oI�/�b�^�_z����E뱥�ˑ�74Nl�үZ�=[�H�q���^�g�/D��� � ,V�uY��;⻮]^_Gg�I!�kLCC�h��(�lB ��u�Z;���4x���-�n�σ�п(���+�JDg<��L�q�ڑgw�Ǜf��z:P�_*�fĔPK����=�	�J��>�ڹ?�7����)����<�Й���x>VH��DQ�U'׿h�Q<��3n�8S��
Nb�ͣ1���0R�u��v���ޭҌNߜ�/���C�&IXs�6����P+��81,������Ƅ��g\ �T�Kx�.����R%�m�ѹ�E���a�f
}�i��c3D����@��:���P��GNF~����S�\�xs9�Ŷ��#G��#1�A�{.��5-�U)F~_(� �6��g�b9;]����L G-PP5�<OW9/7��<g1)�a�ɗG���?+���Қ/���~�ګkLc/��ڝ9G����lm�^�`��-�A�D���v�}$ʘ�>�O��D
-�:��g1�'e��ƥ�����	)]#.��4sX.~��\��^0Nei7�7�<u=a&���Ϫ���K��!QP��=B�.���Ԡ|o�*���ћXt�\�I�㘫-�t<$Ǽ�4��E�G��J�QL���{��3�봰(6V�ߧ�!�i����^_�GYd&N89u ����B@�4�>.�n�ab__�q�>��."�r.B
X�o����FXٱn0@U�*����!���+��ō9蝸 �X��eGHB�$@��n�c�6���}���<5�= VT.���8쑮A�ύ���e)~���L�y��^����)N6�<&ї�B��� �;�<��PfBڏ�)�+�y�)�x`��~�(^�~a��gq�5��Gg|5�ĵ�|��ː��7��+9Zٳ".WV���f[	,�u|Ѭj^�Z����˻��{Bi:�~ޞA�~�aI�h�(�U�R�a��4�'�_�y��	|�)�m��eA�4���\>ZFiu�=B���6�. ��_Τ��A��O꩛bj��?��[�}�z�,;I����XrD���q0�v]N�T��O���/?�+w/9Z�����a��3c������px���V�(t�D�EcS���2s�!Z�)��q MP<_ߍ�M��NdۊSWFMR�Li����{��]�G( ������ȟ)�ɵp�G��Z��Z�J���Li$����ک=Ү%��,sG�F�C5�U��?������:���~�c���1l��������M���W=��N.���E����X��)��u�H/���u�I׭�S8�f���Զ�q����P�A�յ4R�;R=���8��'��E�&����v�qv�q�=�����H9ΩmL_$� ���)s�;���0;�n�z�p�&�_S�J�ج�]T�Ax��%��Rnɑ��yY�/p�G�����Sdm�|�a�����I\��iW7'��l��5?�)�Ŋ9i�	ĝ�e�P���(�|�iYǼ������cy������{�
��-�Db��y30�g�9��Q��@�$#�L��;�)���:e�TK���`?^��
o��I�1#0ɚ�}@����cvp���R����,2[4�Mr����4r�$��`D��u��j=��ӽ'Zމw!ts���JF�4G~�{��x��p�>
0$8�?2|D^|F9b����.��*$ܗJou5�?���*۬X��C|�|�βa��qۖ�ɰL���%#-wpB����N_�v7�/���e�ԹH���kx��]��2��"�D&ܪ�����\�P !y�K'N��:����f��N���$�H��J �?r!�g{�a��b��	���[�2�h�Wg_�c>�i�������A��������-}���]����]*9N�T�n�ť�@c���n��!A�4qM{��y-�q��"�YS�.A����K��""o+hTbC��c�	|��UY�w�GfPK��{��&%w-#Į��u�����ң�l'gn����rD۽+^�ժ����&�A���Ľ4e^�"/��SXμ�
7�_)�l�%?�,�@_�UR�ߙ���$ϴˑ� �a<P?Kۅ�ms�/�4�����l� 
+	h����b̥�����,�J�4�O�r��h F%hX�KZ��`4�ǫ�����n�q��s���@�z3��_���t���z�tf-[l�p��<���eg���5���9#����iG�0;_=� �Nð����,��r��DJʎr������w����:g���@
�>��8�T-�1\D��\y��B
��ɗ�v�*��w���h�:E��	kZ$�5:ҫ���NЏ��J���7p�[Z�>�aBj?5���dA��u��񲻤��Q���ƹzz霒�t�<XlxVHYEB    bf14     c60a�vc}6+"���s��Ci��͂��q�Ś���H�Q�6�z�d�P�VP�%�;��� �ߒ�1^�ܽ^�@�>Ⱦ-1!{xR�k��𪶙R�䴊�-�6_���H��r�b[�����Q%��?�w�^�TБ@P�l�g?lY��n�-|���"S%i�7k`T�1H���眤�[�8P\2��5���L@��ˀ''}�� @��v��Wh��4A�pD.��-_�X����d&�e���)�N�& ��@��6	�S{�J���MCw&�3��+�b��Qz��)4ո���w״���X� Y�]�Ei��xS� �V���6�镓�s��m� �S��4���=!ŉi/�P��A�{�PO�i���t��!��{r�-�Y6p,���G.�oX	��%/ ��t�\�����[_(�{'�K�'�E�mN{��L-��%`��p+�a#���1�4@�_�Ot�� �jp�K[�4e0_���(�#hr�����@���7r��:=) 'J(ݶ(l;��l>�u�"u�-ө�#9`g��O'��&d]+��[���kR���J���?K��W�0�ğ:�-p��EDܣ�)�i��H���t����s�LZ�5�:�	m�d�����q��xf��%�����n$t	U��l<�ȴ���_��dBIB	�OJ]��n��99�Xo�-���rl� ���'͡HM��1�C'�����Ă o��E����76�	�����8h����Ǧ\��}+_z�K�S���4g
]×�#w�XS�ގ{� A��r,��>����E1�Tg�f2�"�K�V��'�r�NkP繳���w��n�V=.��� z2��
���ԅ�f�URn'	0HZ���4�4���=��`�3�>�I�A&O1<�ut<1�7���ߴgW�5��t��32Y�4;�_y�E�e ����p��@*��xb��V�ǘ���|F�� ��m*���ξ�����X�]W��-��e�`+#뎦z��v��k�`��s�7E���7[x�Y������Y���T�-�:
�JL�VՈ2���-%�%�A*g����2����"���ub|�M ����@�0���������N]�r��]�:y��_tQ�,��	琵�~�l\oi�ϕ:/������zڙ��=��38h�	ӡM�k�[?n'��a�	MO]X�����^L�������e!�����A��9���7_3�#����;�I��E�<=�C�`R���Ҧ���j�J�*�װ�����r|*�{�ơ�xu�/^p���ptK\Fs:_�����A;���ۖ�����?c�Ē-B}V� ��aDL�b�KvJ�Lh'����M�-��t5z�.��~$3b�����Y�T�/�c�Y������H8�et:�Bu��AD�ƽ�4�E���/�Ꮗg���=g�}�@@��+n>�.}��F�g��r9�VQcV,a����n�F���T�	輣��HU�U���`��`�c�",:gG�/H%�%�`o$�����D�gA�ڒL�J�Z:=%�ҷ�����g^���p�"���P��{��g��U`:���q�gl	���!d��q��}�Vu��O��)����y<nF�H�d&���6�ǌٳB���j9S�}�dui�}�m�l��Ά����&Zq�=�-|������J�j�sM-�\H<b��&֬r���ȴ�sB�9q�����T���zѦ?'�1%a�x�R�z����o�-Y�V���)��E-@Z��2�2�/m�/�r��*�y�GĩK,8"�&,���6�_6���H9ط
4+�incό�!9��v�U>恾ۊ�~Hn���L~-ќ��/۫��7�=x0��楰��5?��ؿ���ڈ�{Ї+/CvY��1Y��W�?�Q����M�[@���3}�Bo���=��al��5�y������uZ�q:VKg9�� ��+HV�_��|C�^̪U�)k>��?��~�*���hmX�u��Y4��ġy���x�+��QaJ�^mk%��*���&�����e_�|MI�����=��S�X%>sIg@΍�fpn%��}�!e K�˪x��{K_Χ�Lx/a��E�3����?�@�q�y��Z�\s?���ՓGR6%�8�m$wP;t���)s�>l&��T:�ľ�k|�SE�e�gK�������%�����W� _�nsM���,�l˨�H��M�Pd����+� ���y�k�T��r�l˾w��{�I�Z�AU��!�t	��Þƙ�mi&���~�_O����!���ܓс�D�&bB��Υ��U��t����M�����K4�	)q&I\�#\Jy�e�Py� ��!T�?����j^�EL�,�zs��t�Y5���g5� ����3��0�ڜFY��{m��nu�<��W�	��K�uv4gLUÉ����L��&U3�<4��d����j �Oȹ#ջmǞ�]m��93͜S�nG_�������˴(���~\�C�I.�%�~���^���,�|t�s��F���ZF �4ݣ��5ˈ;Aw�+���J�n�I Q��\���b;kb�Q ��I�7�C�ü�kƉ+���AEt��g����ӗ��ڑl��J�/w[Zy<( A��qS��v���,Ց�r�|=�#2k��[ߙ����RW)�+�g�q�_zp0ĥ-z-�XT����m�m��A�1�2Q�sT����1�?{N�|��=ƮP���0��nQ��?�J����z�p9�ῼ+�O3ͱKЮ���S}=E��
,W�%���Te�ZU�\z�R�br��}neӥ�������UlF��x04�K�l�/Q��yxtTs���X||���$(���7ٖG>�6qe�bG�� ��.�2��x?)�ĸ�4�^�EHOт���K.W�e��f�q�h�wB��$����W�Ʊ�ȗ�YU Q�:�o���q���i��y���S9�+]ǘg�ӭf�I�9SF�Eݻ-�nR�$Siw���o�d<g��o���
�ZH|%M--+�a���)Λ��
���f���3�z%�|)���p�!n�L��ϋ��y�!���J¿��-*ր���qT�yW73�$��~q������;��