XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+�@)���:�O�Iv:�a�R��i���;,�`U���fV��k��!i�u���3ᚈ��W����/��^yE�g8�cA��
y:͂�m����"�$^���/�����)���g�W�C��Zg�G��}��5�S�U�6�)L�����g�cケln��a����,�sp��5���7�A��3��ZQ-J�o�=bl�= �������@e��lV3�-1�y�S��M ���8h��WcP0-Z�&OojS���U��7d��=*uփ�tF\���z~�U�C�Ut��I#HOD���{�o��Ux2"��G���o�wV�$<-���Xqn5Jtj��_�D!��1�Kj��&	��Ե� _��i�{?��i�,�q�2~�ꌼf4S�mH`g��xt9�z!��;L$�/Nl|3�v[�*��aK�o8�N���T>���^�]���
���
1�u�=%�в~�(�iP�te������S�C�%�7�L�H�C��n���&.Z0�GN��V8M.\U)��>�I�h�LUŒ����]��x���u�
<��h�y����*�6x�S�(K�N�(�j�j7��7��_������v3t��O�Sg�oV��&�2_bհߦ);�jk4��3�xg�d�T2�0�mf�UH�IE�N��e�9���!Κ�Bwr�~�� C�c�&�����ե	�ߚp'�s@����<J,�u�u���ս���2g��u����p_Td�l�3$�s�5e״`=XlxVHYEB    ea93    1880���idƁ��a!	p)�j��W�&�4E��ŵ�{+��T�2�%%���-��Ҭ�u�HY��	��g�V�[U<�٩��%D���LH�$�I�1UJ�,��' ���iS�fP���c��3߯4<�����?��J��dB���7��;�Ÿ�����HX��dfV�5sw�`�t)���Uք�4�>f��U��.'��u7��8 �N�
����2��"D�E�&$�WIYY@�,�(n۠�#�@p���Yٹ	����2G�7��b����wb�o?�&O���Ϧ�A1��u-��=M�0�6h��(j@�h��[�&��%y������=f��%: �]�����lf�u%.Z~Gl��5z����T|���|�O�|���ƨ��no������ޘ�}�OUS�}�t�Jձ|6��yM;@���e�w��8���� h(��JB>mW�e���'|��z������B�H��-ZLQc��6"kH��%�F����U����"-f��v�M��i��Y��_���=,D���'��d�ݢ�<W�@���3�����7mta�?mU<�|Q�7��ŧŚ���C*'�Pp�7����&�l�F���GC϶�S�t�B&r��z�����ng �ĐX�C�j�l��ْ9{� ��g����!M�[�R����Y����؉*?\��|��At�K��E�Wg�ʳ���P�)UT��FP��^���?L�JA$��5��CK�84>#4�^˷]̣����\I�Y =D���͛ͼ0��S�M�����s�Π�8�+�΋�ӭ_�"�����D[�j�|�t ���$S����~E�"fD׫";��b��>�}�G%��rN>�E���+7�µ|�u��Q�M#Y=`�}��J{ Cn��^{kj���C��"��D��]v;������3�f�,E������\��>[3F���u�xPy1�� ��Z�qH�K�� ;a��(F�3�7L�50�����/�����D�rJC>vIwP5��`ԔWmDh�u�Љ��q�hz����
*�H��5�Q��J��c{U��[��H#����<��KS�S+g���8x���&2�"��9��P0/����vf�I���|J}Eu@H�18�auuu�QDb17�#H	���m)0�E��"q����(��br�A5&�G(m�Q�5��q�y˥r1���C#�i�)��vh�n�.��^����G_�֩ƴ�����*[���¦�*�C%`a�Z�4�A������kG:�-b�~����S	d5tV=P�.�ǻ,͂)�'J���f�N[�{�Z�v��gf���oY���2��f���ݰ�?�Ylw��3A%N�V���X_gk������n�2I��J0Z�,c���ϵh�9���c�QT��u��s7��~/���.�j�].6��_n��M%\���q���e@fz����c��_CC�[螨��GA��|�N*I�d�n|�P�ol5�{���k��
���څ�ڛ���;S��XV.��y&��Fs�ρn��э�Re�8I	�~$_�1/�I�Ye���if� ��"���E��#^�I���I5³�h��"����`�8�w��� ��O{�+If
��7���������j!��y�]u����%�g�M��Hp���W�kBB������h���vI��{v=0!�u _����Qď blTo�%Ȧ��n�����m����#u�t��-;�	������lu~������F���C�ڷ	�O����O��)2<���`:w��&O�#"_2�F[�A�I��t(}񼬑60�e�rQ���ƻ�3op��g�翅�z�	؜F��� ��}k�a��*�u�9�D��&BQ'�iQ�=L˶���:��׮ި�e����bJ%��P��\1�ȤYw��.X*5��O4�&a�x�V���-. C+-Icv��Vy�/���k�t&S���̜�΂/?�i>Js��O�C=��x�O������)B�x�%j.T��t�?�0~|�'�%�30s,y�>4)1؎�0�L��۹���$����ݕ�U��^L����Ф��ʎ�U:�S'��i���h�����Rh4Ő@�� �i�h�v��A[UhS��@(Sw��</�r]�Y�gPb�X&*V^�Э��h���3Lf^���{���
)��#�R��\���m:�T�I��M�FD-�'0b�y��WKm�o�k�M�{�����H�@<��VZZэ��c������`3^e��L@��3Jz����p���-Q�:Y�K�>��np���`&�5���[k���Lѥ4TjӠ���ެ�e�s2xm�L�_�<���=*ex7��KV��=�|�#Dc�ӊ�^B̈́6���6]�/�6ї���.�j뒫������u�����l����ɧ�nM�H/��S�o�%v����,T`�hk�iN�[t�t�q�'D�g�mق��-9R�Zn�0���L�oR��bfd݊�L�Zv��6�h����"�z����Z�ht�Ǵ���V�~2P?�	B��p��V$z*�HNU����7 F�p]��S}_�Y0�ṭ�餑q}�ڮXPWw��ќ����)I�y���B#�KC�.]�W1��\^2�nu��T+S����
�f��k�b|\�������D�@J���I��G2�䕴kt_�>yN��洷��?��c����.���5�\� �1$��D��!�)���H4�8@���u��ZE?���,g�wb�t��3�V'��8{a�t���9��}|����c�E��B�o�EZ���h�;Sr9Ys�������X�]m��=s�d3� �	 ��A��ٍ�oހ�X¢/�K�=R���WA��u��W��`� �҉�\����������Y������v, !�\��^����Ap\Voྔ7ik�'�0<SG�T��������*�4B�G�:��@����[SMb?&4۠����h�M~�����\��S�{��!��E��z+�|r�ճ�����(�l
$)N�� ��i��K]EnXݚ�Ԅ�<劐��I��_��c�#�"����0&���ϼ�3���$�8�T*��ɰjb��=N N��ȳ}��Mb�C�����H_�jo�[vq��*�Daɪ��(탾�G��N��6	��H:Ʃ���ڻU�H@��SOy��(��ƆK�ֽ|�x9��e��H���/�3SV%��$�e�t��Ε^|n�5y��������Է[�욘�aS~��2��i���Ǡ_��i�לm(�AK��_���p[�Ʋ�V�Al��D5�L��
0F�cIz���#��/f~���W�',�_�q������(M�??V��5�;������/��ay���l��D�zU���"��7^�9ՔO1]�	Io�~ݽj�BB�_���P��d.���v�;�JpDv�iX��m�efHl�p�j4y�͜�=�K�D����w�@�"¥���ήd��u8r�3)��b]�Q�a8��˫[@�߷����;� �2o�m=�JK}8��z^�%'F��f�S��\�^ښ�X�B��I� �R������m����p��2�#��q
��a`��`H�+��zO\J,�5ͥ�Z��Ѕ��	:q�`� <m�r���NWQY��2n�p�0�F��Uo��Y���*���S�bfŕ9���KX�3�������������521>`�s�%n�����W-s��5V+���$�7��Ņo��\��"��$����-�7�?Eo��U�Bs`�,Q P$��SSl����_b>'.t���^��~�X�E	�,�`"F���[���ρ:F��X������	����7�o��9�<��T*�w?*P*b����Oʇ�� e�<��8�t�v�.�S�'�{��P��X1]#{���K����V��ʙ���&+�/E�q�8��� �h#�Wۜn��Tׇ}�V$??�U��H`w��C,E��h�j�Ɖ�Gn���r��kf�x9㏟I^�Vo�з|�����kp��{-� n�1i�s���Y0�>6�'5�'���z����S� I��wY�7/�+Oܰ�P{�t2�I���4)�+d 	���4/�d%����P �5DV�{�TõH��'oa���Yh��7�����qĒ��]	dL�F�Xp3�!�:"��؀�2ZcH1(_5���\?i�')cY�ꥩ^�S�%x,��w�ӈ`���&,���/h���	�@v{3���{���IB䉵C�hi�Tc��}�BizL�h�
�z۹�)I8�
�|�n�+�u�5M 
��He�^ ���*���90�r���� �El@�������g���?�*Y[R��71ˤ沸�� ���ӎL}��%���9�ȅ`N��y���6iI�Bh��z�� f�V�*�W/8���Ҕ�F���4�{�uUo���,��-����!��HB:��a���oѹ���G4�G����l�g\�~[��0���ȶ8<��#�����_�TfW#��Ij)���D�u"����go�qَ���,�̷o�`\醜��M��/΂>�EJuʇ�X`�\5S�^�v/�gzW��n���C&v���S�փ?'@���xw}��\�M/�?���|�q��zgi�RsJQ�[ *�aBٚF+ʤBB2� 1y�j��'�}��':�DW��Ә!�1���A�#�_?�R������~���Z��U�쪼�36����X,���ʹK;���z��mX�}�62��1�B����/)���=
��v�K�9<���C2	�TV����|C��Y�xO�tǝS̂�E��Zv�j��W�">-%����3ȫ8V�ٯ�=̼뎋�	sw$d=��p���J�ao}6����?(�������y����`$-��XAP�p�n0u�t���e��$���)'����:�оHr�<4R��?4)Dt��R���e�7���}���L�y���_%,t�#�@����L���?Y��h�����$B�5-��~^��a:��|���?<?��n�Jc�V�2�@�(�r�_�H��f�9�(�k\���kE�i[+�kt5��O��~R�Xғ���U��T���ةU�f�U4��=����Q�T%-����_��:�y-3�֎G����cݴ7�H6��#WW������I����#z|u����;���ҟ��#4�BQ��o��*�k�`�m����;i�y��7�YW�V����%��7.�50C4�K�JK�h�L@l�F�����\��,D�4��dy��-r��?o'��ft)Rl�p�n���A`�����,y�^�jte� �<��1� ���z4z[7z�v���߄�2S`����l�f�G)�O_5&n��9�� +Cc����u�d\��1�y�O�Ͽ}x�U���K2 ��#����x��/�%�@t�����N���8��p&����Bl:�n���f>��z`����I�L����%e�@�"�P��<��*���}!���P{f��b�O-�_,�&�+u���6ϲCJh�T��5j����e}MT��[d��5eD[��F?;r��P�#�-�a�k�!�vmy�a��R��~�4��� ^��V0	���{/-�ZU/_n��N�дc&p^����`��=Π
!�D�C/�?�2L
�#������.^�ג�	��8�H�%�Ź�>:;��
�=0�q෶��~����ҙ���^����A�!���#6J��о��%�ޜ�P��%�VԃxmY'��#ͪ)#�`���x��Tw��le�������C����ՁD{���y�x��Є��r@�y�����§�"?ı��U{��w�)q��2��6��m�âkG]+�%*v-+h�نP����p�6������Y~��QSB��]�l5��ug�s��D�N�;r����V�?��2��
%ewҕ]�p�z��.)|��Ȇ2��끲�%�[�;Jeޗ�Ɯ�Za�:Q�f�)�C���ATp��j���F6����b�\�wR8��j0��T�� �^Q�,u�2ɏ�Xґh7/�hCN��.p��[W�'�����#Ưy_b���P�E��׿�mzj��e{a}� �jCJR��N�N�Mp�\uS`kؤ�