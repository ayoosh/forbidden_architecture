XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|�9�*6�GN�M���ĸp�h���_�m/���l��M��j�e�#o��=x��=�z�.ۍ����>��x��/|L0����M�_�]�<42��Ԩǜ��B*�P=
�Y}��k)]�7�>�/EN
�,Au��+��S��������8-D'��*Yݜ]�s�~��K�'����U����;��Ɍ�}��p�yxC�����ԳZE�+�PJ���z�Ǥ�/�t2���[_��BŸc���8t�3U�zl0|c⥭:��\�N7!�h?E��sĿ��h�Ţ~?��d֪����g���R�_��s�b-�h0���t7�!�(��`&�gD�8�K��U.N="�<#��O�����0�J(j�92v���_n��V�Ѯؖ]�ޛ�g���*���Im���JĜ�4�V3�&���O0q	vl��z��Y!HP�k�(`�f�6����Q��p�5�JqTj���F9!t��ƍ���pI�I8Qm2R|�F1,0�-�l]�.>o�7XQ?�q�,ϛ̎���Ø���L޲�{��G̑5@ �H���*Q�m@L�5�ȩo�ǰGK(�>����@5|�������N=����������̫����Ư؈�&E�M�	ml�8���|��
�Qk���|�s{$�c�[Z��A���-�*Ss2�2�d& 1DP��v���&�[�_�@6�S�.p�B�Ss�_A��(LOi4#�*m )���b�܎�mгK_H�:M�&zz|�^䓵��)	XlxVHYEB    3504     cb0nh��_�s ��{"�~:IE��f>�v��p�*s�i�}xE�㜫8s��ctC2��!��[O�
��I�]�T�+*m+���-Υ����T�NG�m̯�����Ye(�I(<Kg��q�n�e��B��6F��r�U�/�3����&]�伧1�;�:@[���1i��`�LX�mw�?6*�.a*��Sz�EkNU�n�xe?��ۛ�ӣ����gՍiA�G�nM~��L!� p��9�uj����A���I�3[i.(-}Q��F�����t�M%�0M1��#?�N��G��e�Iu�w@UL.A��
z�ud�[����x�5���@�6���)�
\8׎X�����T��O5KD1�"�r�*�,�@���6[f0\S��x��Uq�a���{9��u���UPۗ�@iw�ziE]�����mK9�%	�L�{���#G:��n¡IР�N��Ĉ6�p�̬�
�J>~R}h�ɇ���(�BkG7v�����@Ⰹ�����;
iY�F
6��s"�����Ǌ?K��2O������U���9ڹ
貉��5G��������:�y`"���UQ��-f,q"�4$�Y��qqVڂ#a\X�~PU:R���/��FdS{/>&��︚�ϗt�z�4X⧺Z/
����՜Q��txC�{������y�4OD�/	��X�(�C�V��~��-@-��hDc�<�D6����#�>B�h�o�����ۈ�+��:P/���V.:r
x|.�"�2DY�Ď�{8�Ĳ�9�Kg�H�2����Jt2�W&O�����P,����0�:SCr)�9�� ��aIC��|U��Gg��TN\E��V��ʞ�\���#d�}B�� }�N�I�-0���բՏ�u\���R͆De��cU����>��(j"��`��2C�e�L-�R��K�&�����S��c�H�����h���=Id�;�w����Ev�u�AAԹ��ɫ�d��;. �k�����N�+q5J�N��~ja�G����Ht�eK�OE���4�%I��ӎ�����cH�C=-HDgƢ#&>�9�k�Vx��Ђ���I�g�t{bb�Q<��?�	���ty3�y.W��(��E�,)�O-g;�����gX�6Z)疑�u֮�,b`T\z~ih@�ԙUf'}���
�U�^�@��D�����ü<�
N&�N�4r�D8���^�¢~�K]��s�:���s�1��z<�rb�{��#���Sl����5ݍ��G��/z%������\���Mf1p�VUC�N}؛)�Z_�l�h5p'~�6��{�����2J_�����,��m�VySUV¡*�h�� �yܙ����B�l���_
�V���6V����� n(K_���R�d�� :�ݾ�5'��8�cU��"��P�e#o�*�X����;nѨ.��4ʕ�������B35h�[pʝ1�6!pW�% ���`��tp/r
���1�����>r�U�GړH	��1>���|3W'�� 9��_�ޮ��/ٿ�6��]7ab��W
����uA����𒆤`Пax"g�Rqc�	��6������_筚���jߦ8�sT-`�F?
�w}^�큊��,�g�CXc�)7I��5jo��(��$1�#MO�F���<��שZn�� *�y�9����6K6��X�Ě�����X�0�-KB�1�
ٶ��ٯ��U,dl2�0]VL����[��B�ʣ�\���$퍦=��8��|>/�+g���]I�w��T�-̎����˱9d�������6������F�Ic�z��K��è���yj���[� +֚�U}��q����k�C">�3mh'ݎ�4�&N_�Zv�ڑ��I����V1�"�I�t���߄ ����n�N��ӡk�Va�H��;���F����82�9��z^rʺ��`-��Dٰ�r�^5v�BU޴�j#�'��w%]��Љ�� Ufȡ�V�F?�qrF���秃��������4�[�o�m@���HF�R����d *�z� �R��=tr��FI��um�<��Cj��n���P��	U]T�V�2T(�b>����iB
ɍ[&@3�$�,�V	a�o�r7�϶"��Z�y��w=q
u4��dG0��E���|�č���K�oٿ��B"kOi��:! ��wS	���0���;��83y`�,<���E8�}wEx�|
4D�9��?{3�
��i8�h��;7�A���7,�
1�W�����8p�/7���N�ﾴ���d&�����6�J����WϠg�u(�]FP9����d���+>�i����Z��N�w N�Ӆ�酼�?e�f2�5X��i"�4A��v߁U���x�.+�:EY����˃�
AM�4�R��_7g�)9��4U�ْ[��w�t����4܍JR��%�"�{�ˠ��2+����<*敜|�����:Ԇ�
ֆ�P�`�V�}�>�, �\+�(��s���j���P#.P`cS��Nv�T<�G8�N��	������QVF9a�*�#���ǀ���3�!���oX̆d�/�B�MO������l^����bF%����,*%��_�b"����KM�=�[�U�(*���]����24:0�6�L��zG֜k?:N�*�_ğ��bR~f�����-���x�mC|�����/
_��վ�׻q��q衛�j5�D"+!ya c��4��@���`�]#�g5�Ȕ�W�]8MS��aĎ��
H���pyNҭ{��xˁ�M�)�:�^;_;���T�?��ХR�d4�Bɍ|��-Eh�8ɍ��Y�)ݓ#R�	X��w�ZgjW4�{��s�G��J����LK-x�o2�c(7��E��s12IR�2ǀ�,]E��- �o�~�`L<~�.�,�{�
��/�$q�N�����=��`�bS,;�p�qD�,\桟B/��Yr�S�1۷Du+�ֈ6�#�[!\�S�ҙ����`��6������d>}P�f�t-HOc�E�08I1Zj�|ds����32�hd�I�+4�tT��|3[�!'qnA(�Z��(�e�B��
xR]�F��{�O�{����Mj�fBh��=�;(�\�U��4�^�m<N��7�*��|����VqS��'M!ϯ�r�����E\d��Q�_��?j ���o�#����Ave�l9<+�1�l|wF�{�B�