XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��UnݖoV�|�ZIȱ�b���\��㡬��U�(H�C�0J���/��s6k2�>��H�o��ݑ(~@C&�E��0�j�7_����y��p��r��!� �'�X]I�S�~�h���VK�*�K;�
��v�V�����3c�Ӛ�<I�pm��(FT�8T]U����ºm�3�&ۓ�z����:��S�����ݢ�el k�[zf������J/qF�� c`���]k�w�	�c�(�P�$1g�N�*Z	ٗN��+�iA�#�N4��^��l��A�|�zN�+�V�=�je�A�����-yz��\��W'��S�_7�IP7DQ�Z.G5��6�u�橀N彪�+�QZ�_tRb�Tc>l��<>�IM�
�NOV?�R�(_g����o�8α��0(�c��/����>���ER�3��Siƭ']�� ���˴A�)z�pR�k6�hx-D��np�0w�W6>���K.@�¸~�g��NW�D����Q��]4�������JD��mc��$P+9)��J�?;H�s^�C��&?Zr��+g5�P�J-�y�!_k��\m��u��!����V��̴;p���v�m�G�C�c�zC��7���R�\7�%���JK��_ŉ��l�0ʿ�����|X�D%A�I��������B
ir�~���>h�QQi��N��]�'�e�y��f'[��Aʏ�AZ�|�I�=[��Ʊ���m�o�׿q�jA]�.$-�&L>��.�[G��R�&�I�Eڨ����XlxVHYEB    b8bb    1ad0����<F�r��2�kezu>�nu>|�4����Xm�5͑fh��B	������m�t�4O���2�����KEJ�*�53�LvX�_�<�^lc$Ѳ�q�� �f�\���Ғ�B�M��U�ܮ��3�/��		c��8���
�|�K��P�/dZC�I���A|���"̩W�,`���&��@d&��`�����_-�f�����k%���N���ȂϷTl��o��:w���<��5�TL����A�t���99�AD�vX�G#����;hW���[�jPX�t�j�O�#:���Y
~=;��j�N��l�,2&�<^9���H�+�Ғ:����k���Kp�Dئ�����"����ndh�r"^���z}�� ���==����B�oW�]���ih�}��D���N�����vqs��	������8�� ?��P�Cj)v	,��Q7��c�?�e�D^j�\��+Q��hܥ�"4k�~�B]>���]O���sF�� ��o��D� | �:WXT8�c4m��\���V�J�HI��C��]��=��⋅j���k�T�����5��c����c�e+*�K%/KD0�vs���b�
A+AA��S��|��a����I���鳪�ޭ3������A����y�wG�A9��hj�!�*��f��=��bc����=�;��������q�!F�5���׀�	��m��a��.������GûL�c��v�$?ZgQ����&:Ū�5�&����ե2��Ex{�Ӌ��|�W	��H���Fw|(�ȧ����+� l�(j���W�1�e�����:���83��/�sU���X���������S8領nkݣE'�F�d�?��o	��r�;@�J�[]�ɩ�f��<��8�VL�40Xu��IMM:�OO��p����3����G��5,�Y�[yS�{��ET-*�o:�t�#�	�+O��:��K��'��93�~�|�p��x�<��)e�a(�"��qė�d�rQ�f����x�q�̽9�m§Xm�S��a@i!sw�����uT5Zz��_c��8)O񏢰����.uu�=Q�~nT�o�Ґ�9%Ok�����:{B���0��_���A�����l�S�ܤ��o��YG� ^,�W�y���	�s��r� EZ�-#����v�b('yb�`a6]i-�3��DKr��;��X|��5�E�����6+�mS�0��]-��8��)��蹁�k��f`O#6�䡮F�T�/���W�Ň�#��0��M����a�e2�Fpu|�L�Q�-��gJ�_��r&h}�J�MM_��+�q�����Pd��(�Ѧ��,r�p}��f5�[��N.g'���[��|+���:\�ds�7!�24�"��'�0��� �x˂e�$�2���}�����Dŗ��z��2oQ�6%G?���/��"�����i+v��q��}��No�X��\��G�@�Ej>�|By�h�8Atf���&y��#I����U<P�M�}���m%��g���3���[���,�^XF����9e�(���uH�G��z�˂Mp����������]���,Y�Ԝ]f"9�i�/�@vhF�a���	���B@�(��?�_5�G2Z���Q®�=�8Z������`�Jlؘ~�M��t�� ):m��4���w#���v�]�S/̲�~�q� ��?2T�<LN���v�;�:�-E��z��vy?�:�)T���p�|�u���V�v����~�J}PvKKG:��- ��ތ�U:�l��_{��$��s]�ˈ�&��=I�o��؝��a8ܮۅ�m��sٌ6��E~DIp�$ C��f�K�;�U�����Ӝӗ�����GS��������������r���0t�R�~�O��a��g�,��.P����p�C#@��l��l������HHP�)����R�Eɔ�x����k����:mX��2���?0�������s��e����C�)"�]� ���j}�h4�?k�G<���m�D_�(���+粅�)���t:�H�~D��	}�BP��_A7�so���M��2��n��s�b�.�~:C:-#�18���A��e��m��J��0�D�Q��@R��&?��h�˲�����P`�9	�@�^��7XIjZU���= 0��T�Q��x� �_�HM#���A��Q��׊6��52���kg����>�S2X�
%e)��5�3�<}�
�U�O(�V�Dc���Lkz�k�};�FI��֐�0̃&�)�:X�حJ��?�v'�T�|;�<a���n;�~6��x/oEk`"h�R5`�B�P�@�48&C��0�C�#�ء����"{�p����꾣�Z#���@�i$� �U�h-�B�_j��ތ���#πP�C�+1w�V�z�&KƏ ��L~��q폅E.Ƶ�,�ɮ���aT%ۦ=�VM��{��G@d��d�m6�-f���<�Oy�ߒ��^qG����'Wy(˕�~�^\[�#X�F�l�/���Cj�#֣J_��\��n��r��,f�К��q���wo	�i��=9x�hɳX<���R�Ǌ��*ulщ�><����(����tW�Y'����[�z�{���?ja-R(0��.e����'�+Mg���`*�(C�ґHUX2�ǘ��ٱi�,QKF�#��&#��b��TX��Ļ:�
��W���`b���ղ%�8H��d�=��\���e�����e�F@�5�)6�ƿU�q�o�nw�:!NN��_��\]Aq,ݳP d��o�	���ld����9!B��\;��{{�B#5
��FwyS�B�9���0�0�wT��=y˅Ԝ����;7��U�R�w@���H�����zjᔹ2����	��?�[&ֹM��f'+,B�����euG�#��#���!_s0}����2�����=�a^���o�C������~<���zچ��C/2�l?�sX�@B5cQ`Kh���n��a؛/��`Ws	�I 7���^�����P_n�}�*/oq�K1�e�.�S�q��18?Vҍ���#�Sǅ'm�W]Ĕ����w�{� <&1^
�>�Z�K!��� ��)< 檒���2sI���oҋk\,X���Y#���<~��ڏGN��[N���(�E�i&�xL`�gO	LJٝ�.�����D�-�Ơ�A-��p{��|_ȡ����Mk86�|:��>�b11b��q���/��m2����qҰU���zu����� ���D�W��_�)�T-�d����6�k�qB>"��4���z���JX����>�)S�ȱ(��9�Ů��'	ǓJK�����M`ǔ6u��ϻz��c̟��2ԋ��~ƚ�ϗ/���
"0�;�~@h�8X|<Wؗ�Q*�]��	ƛ�j7�F��c�FD��H7��	�<o�,���
��>���p�Ϋ�f��t����`�V���V{�Ę#��T��-��ʇFSg�L�}�K֒��K�LA9��Fd#���mLn��Ď�}i����R�U-���S��%��J>���|� �m���yMz������ސ��&��<�`�S#\<�=�� �JpҀ�Zi�:�{�S^��b+fu�����b������I����_T����������z���Gʀ^���^N���8��bOFr�֥0��¨�,�x�t����۲�$��[���EVu%͗uͼ�We��v,�������Ǹ��i�_zS`~��}p ]L�|�b�!��UW���d�&�r$�"��!��1��nǺ��AB����7즁@��k�0���&F߰Q��=���e2*�2�,*v8���n~�1<K0a>����\�X�7��a7g���2ԛ8=��n�8yʏ$��F{���N�hT�%2m�:>�"�>�
��=YX�h����ݧݍv�R�t���um�3��ݭy��P�]8[ )0���7�xk�2L���a��̃<���wl�����;��)�%K�#���9s\�X��q��E��}�����A{aO* �e5*B:Z-gd�n�����ŗ�u܃T*`�B��뤽�B
�n*u���W	���F"��YY�?+Nӿ{��ffͻGں���v��������Q�G��ai|�	�{}�����.P�LR�Z��x|��u�`{q4�$1X#�`[[�t6)q�;��c?M��Q8�8׆؎iv%Z�a�^-�!@���=UF�H�4�뮒���k�7�a��[!��ݥ�<\x�W"�j9S��ۍT�Μ��4�?9 Th�U^GR|h7��@��$�bT6%AD6ِ.|s�%�_R������O([ݘ��-Xت�I�0�nCǗ�L�5��ZI�}��j9$���c��ms�5��rH�S�N�a����Y�(�Wl溏ԺF;h7�
M?��-3C�O���\�a���8	��*}�h��`�LE88լU�bFE>S�Mz���pu#�\�#����I9�{6�.)��0)됆�'w��sįt~qF#b�����m�n�ߨ���C�ȯ�\�cؘ��W��Y������	�TS������P�I��ݍ<� 1��+����F�O�~Y�$(0G��"Q�73 �Ũ���w��R�ӟf�����?b.�#O/�D�9=�����m�?��LX��RxhZwI}�^���� .�����n8,�Q=x�5�%-�m�9y@k�a���glm�W�-�N���B.�%pu��4B�3	>}őS�<�@(�oQ$�j����j�eay�t�Z�H��{��B܉�;[b=b��prn5��bq"�\D�f�)+�BN�^��(b��C#���U��3�o�}nZ���$CE��~e2��+.~�c�L'�t��%ҩX6@ZaV\k3h�}8�6�ᅟ	qJ���C	*���RS�M����h.s ��9#d�V�s䝪dǾ�T��$ 6�᳛J��>�ҟ?u�]]�EՃ��c�	B銄Q�q��-�촼��@�I�R�'�6va-��q�yWQH5�~�����7f@��.��0�������i��4K�]��?��h+�rzC��$X��pCugdX�� ��o��+��c�y#���C�Ӕ���Ӷ�2Qo��+;���&�R/��6�Ө�8�&j�f�݌X!a\#p�f�ߢ�@P���:��s��o38�-��l'伙טM�6�h�T2./�6IL�{^�_��~$#���jtd�ڥmd}� b��f=LDd=�l�"%��OV8G��Io	�m�����������8��V<CJ�k��v�L���:��0C%�P�4�Q?x�^�=N�(X����r /�]��=��]M�8��bJ��]dVt��<e��^��ےV��\�lI>��~]���Ő#/�U��!S�Y���v�ҹ޽��b_z�Zi��M�5�}��c�X�ST2�X��9�\�>S:.Gb�pX`�R��y'��%}�C�Y��yװe)r���B�ZN��Om��ͫfc�tT���4, ���ۗ�~�
#��bY	#	Û�#PG��m��v|n@�X�u2�y���ݫā����̛���:s�~�3�� 0!��o|D��̙��.�:�d�������cއ�[_�dx�S�_]EU�a��K�+�����Ϩ���25E���ʯoFN>_�6j�<�ǚG=a����ضC.��$��Dܡ�͹�d��>��O��aW������n�"!����&��|;jө1>�=Ы�W���R�IW�o�M��u)N�b1~�F��Z�����
̕��2�
>�;�`�&�=O�[��@�����3;f!��<�D��=�"��M�`�{Mr�=Ñ-��[.�.�n���í���7������))a�|���2�M��!���5�=I/ux�J��� Χͥ�B�*
$��ݹ4	J.��<	�}�}�Y���ZN_������gT���=�_I/�r�'�W�)ݮk#>4���r4�!� �����:�`�~,�(~�u�N�<v�v�+�k)������۸��H{ �~:�����ǯ��bOlYv��#'�����%i���<�z5XK�´��g�X*йmr� �cTg8][Ѳ&I����:xՔV[BH���b�D.T��Y�F�!�s`�nŢ<�|ű�
�9w��~$>p�R�0�>w�EeI��LV[~�^P���ɫ���b��`�LmN�����<w`:�?��I�ך��DS�л�(<2�[͙�%j�G��C�u�/���[h�����j�l��X���l#�Ů��W�|M���)�a���\\����k��#޼��0s\�f��gK��]R������8.ѿ�`F�J)�0��CN,TY6�w�����7t�sВ�G�����x{��e-B(c��	�����c�/l8��ܳ��=A���$�7�7�~�mJ��Ւ<֭Ӊa)^u���˷(����۬�d�s�:��]���0�(�Q��k����Ch�4[m���)t��r?ǔ������+�!�Fj�.s��ɉW�~�j��y��#N7韲�׹���:G��hu������]���e��¬������$���l�M�$N��"�5�r��ZWrfn!��b[�.�����2�h����g�D���x�
:�Q�7[���[��=��x>��2|����v'"JJ"��P����w�aT��rq�k1��|h|�0�i�������