XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����֩X�"j:���,���Ct�ו]C�k(%ab�zU�������e���M٧��P$x3W��o�K�������{��QF��G�a��z1|��=��)[Zu<���Z3�����E�Zޕ� I/r�`�\n�-�&#5��˟ї_b\)��M�/E�!���z���D��r�����5F��$����J�"�ѻ"�{�*�N)l�(�?��k�+g�YjUK�hmL4���!<��#R�iuml����r Ck�T ����p^|5
�f�>ye&�0��G�b��&����m�{�)c4*��4�:9���$M9�&�f��?� �C��r�X܊�jN0<b���z�u=+R��D#Ƨ?/P�E�kt�;����bZ3}h,2�N�g�(=BK%1��B!��W����R�$%�4<Y�=f\S
D-f��/�-ܾ&0�B�~��Y����|L��J�\�ک��]���O�64���u�B�D߶qͿ�Dst�N����fh�2-�!������:����m��ӁIX|�iq{Z&�����Ȭn�&�	A3���$�.�t�m��XoA�]mW�-�4W�r��Ǥ�Z�;732���v�3���s9�;�6,۰����N-\������3g肂-6�ԅ�3��w\�Z�l��rֻ���3{�Rr�5�=e����s��D'������d���'M��M��k��.�w>:�2z�6�BX!��l�/Q���˚�H/dk=٢DQ}0
.��!lQ���I1&�;G�!(݀XlxVHYEB    fa00    2910�uB�y�;�aA�=����Gv�ղ�����L0���nx����MF���(�	��Q�]���0Pl����`ӽQY]��ܩ{e�珰���}$}���ǩP1~���~Dݥ���>&�i���O�^j�G;��i� q�	����h_|*N�=ۙ���=pD�b4,��k�L�����T�]�0��֠@s�k�@׌>�/'j�TF"�ȃCǡ|�mJ�����*��>����B��6Bb��$�j栅^G�58B�w# 7�.I�0C�2��$�SdJ�M�S!~�0p�D��|8���6:��0L�q:�{��R�&sk;��}�h޸�1-��(�wC�lא���/Eqf���������(�)Q2j��`���U0y�v�w&�U��1r�F%��_IzBu����'S�S����2"~Jhn� �F�@������:�d���&��v�$�H����D���@�6�0T�V	��2q^p��Q�.��4Dl�����{����XJ�Vf����*���#\���v���8�
ߑo��B3f~k���AJ4�R�N%po� ���Q���USgB$�f�h!F`7#��C�[������]�����4z�����Ue�n~��MghŊMp
lwI߱�����e���v�1�$9�}̟Kn�@�˙��A.����}]h�<�c�EA�w�`eTn�F�QL����Z�����q�,��?�1���lΈ�6%~��s|}�$
�.sT֨pݮ'Ȧ����1���U��~��U�Q�&�m8�4��f���!,��+��S��2pMdy��@�	k������l��{Z�~$.��e�� hs)M:m(*�|z�}̳����ٜʹe:NB��eԹ2r��N��n�Z�8�&D�5ȁd��k� խ��p`��k!�l�*��	 w$vG��9�%�pA^��Ud�, hV5~�W�3;X��u[�'�"�@;P%C8	��|la7<c7�B�Ȑ;�_8���"\��"+T����� ��|�DB���L�x�3�����Y���$7M_��	�m$.��Kz��L^��\�jA�^���Hew����&6t��lv�g'R��L�+�tROg�~fD0��M�H��0s=�4�F�� ���D�^�]p��E��h�RA(b��g��Q��xo��N9��p�k� l2m�d���U�=�^I��"���~ȝg���n��|.
�����IMi�f��?P�di��og�Hzi!V\��0�2XY}6�/E��2�(�E��3�r��)�L��z����Kn�*�e��e@�H^ _�]���ဩ����xr3�Ճ �����,ǌ�����k@�W�l*�112�L��-�uŝD?��D�ͷ5����w�U�2�����)N���\wᐖ`�`VUg�x�b�l�p6��L����H�3���Y��� 0�(m�EC�i�y� W�Ow[�.��d]��<2��5Q�4�|&&��ڄ5�a�M�6!ᥕn�Q��]�Vi�"�x�*,�
��(z����/Λ����e�]�3n����&L��0�Ix�;����YP�K�ܒl����R�
�M�W�d�m�n���A]� ��Lu�S|���tБ� e��������R��9��9�ށu΢�b�,(1u+�]dNt}f��Rl�t�	�Cu<��_&\u@.ؘj0�* �@�����(�_6���j��3�%��e���qߥ�y�)�A�4d�}�N��b���<pO�E��O"���0�Џ�e�&�*gl�Lp�dh+׳�}�=Nt���6	é�UD�����@��%�]��� ��2��/ �pZV_�m^��Ѥu]F2��Ả����X�����A��s�]��rr��܉(j�x��H�; -"ߚ�+��uD &�}��n�V�Bd�c�&�#5�߅6�[6���*���N-;#��}��f&w_�'A�K��:���%:&A��䵝�A�Ѡ�ʬqm����h�L	t�O�%s�!�n�ZW��9Ԍ]���x�h (��̕���S�Wճ�}dp�hv�=���.X�5�9 Ӑsj�"~/^�X�_4�<�h~ j4h�u��w��מ�&�,m��U]=��	�"f׈�"��*S(|���B��!`3GjyV��gre_�l�֞�W�W�,(/�c�R���e
�{w�}���W̗E+�	�w6���c�s���@���6�JnL�6�N�ItoV�s�6"�rD��X,��@�C��������k1L�G����|<�Qj�
�r�X[��&]n��. ��ai;�V�)Ț$g�"�UDȜ�mf�$�y��UC��u�
�1K ;��reR~Sٌ�S��}��#��f���6O��GnMx�m8,(U4����q�?��cI�n�$���Bя����"��(zo�V�1k��7<Ƣ\f�vg �50���T)�����e�Y}��z`�;���n�.4���s��s����Έ���,�A�c�I�ɍ Xd��:́`嫅ƌl���Nq�����@�Os{�IJO�N����JH��|���/7.��Hj_�>?����1U1d����:&%��$>Zo��t���=G��Iz
�RH��#
����������ZB�U �������3��`1�����B�4��4�"}��D�a3�B��H/�H='h4�f�{�r�byQl�#��<���'R��V��Z�T��g��s-���r냔�5�6iYwaX�EQ����u�a,�O�@p�����x��/�I���um�]	c�o�'����i�~,iEpA{��n�L���m��j"�� �j��C6Y����8��9���U��U��w?mK�k7T<c�VC�k�H꿻
���-�ٱ�*���ЃI��u&�׼��_n,Y{V
l��S����7��pn��w����ɪ�ķF�{����e�Ā�T�JO�hY��R�i��X���b���u(��/�@��M!J)�΄�H��˚)ګ^C�[�M�*�o���?��ǆ��ܮ�������F��E5�ղ�\R���<���8AF����.�=U�E��&�Hf����9m$��1��r�ce_�kKZ����,t�R���Qi݌D� ?5{���[�Ŕ�HoͶ�ݾz�loh�6�j�e���B���C(TdC�(.D�x�h3z��-!�88������+~��Sg�_:�֌D7sGq1��?�󲨚{fD��'	_p���'6���L����tY�h�I�C��<����4��=je�=��~���p�eK�S7�Nm����T�E�V�m�h/��b� �	�o5ˍ� �G��(\���ё>�w�2$]�x��M��_���o C٩A�>������]Q��M�\+j���&Z_Yn�����/-`�bnf	6��%�S\�j(���,�/*m��=	�>ə�4��ެ=|�0���ڶi��y�*��t�L�%�ܓ�J���Z��l1+�і�Wue���(��S�:�V���ogO�Ohq1�<X�R�����:q�,z��@l��O2�����gjߏ��ٍ
��o����V����*Eq3�P$�[�R��>�.Sj'�x����΀��I�Sϴ5�����z����3��%~�n���-�F�C����:#i���C\��'姑� �<���m1݁��}aU��!9Y��&�TMN��үp��n^��p75L�K�+�i����*�lύfos-�5BT��1G�;�@&׬��w��0�<3S4b���UP$K{8M�xP�x!���Bw����Ѱ2"�-e����<6֕l#�5�E�YU�3a1(̥�r�7'�o$���+3�7lXMۥʷ�l�{�E[���͡��z�&��,-�}�ZVR�sĜ�������r��[�x(����m�g�:�R�����w�)�L}B��8Kٱ�}��S.��L�3yxcGy�����W����H�{C��0���7j�I�C�����w��W�z�+�[҂����d�]�����DƕE먺Q#���܃RK6];v�0p{�f]��-��;�p�p��i0��v�X"f�˿r�7����\&#��!�ޒ!) /���<hD�&���ì2�)�3E���kG��Êbܾ6�f�����T�����Y�`�΃qpU��so]�]�0|`&�cY���#���i�XͰk^LɌX(7hO�la .k"^�.�U��ko��8E��M�9�b��ʂ�x�r��,,�6e���kޡ4p[9g2 �!]{��t�W>e�{��&�ͫKP{Q|ò$�t��t��m��s��y��7�L���uO��I��:���^Fg�R"I�쩉)���=)���;�E'��nP�����P�9ٜSȻ�Ʊ^{�s/ş��H	�sK�p��y�WXtbceRK%d�5��$���:�7�Y�+��6�B<��b��+���Y�Q]����#�m��x��
���Y�Ɣ<g�c��/e���m�O��t̓������{�X�c�B�|D6���X=-�jW81�J���,��pMx{y����Mq�{��pܼR9ɁR�d��� ��p�{ㄵU�x4�G}�c��1!Bi��V�F�ى�y��k� ����\�c�n�}�9�JP$�EK�@,��B
2%�ˁ�+����s�V�(\�Y�^.�@�8�W���g����2��5���Kzz�G�5�����P�tvD�:�[� {Ea�="�'�c�A��o�٘S�C�d�To�O������ݜ��;[;���LeQ��Z�U��M�s�L�mR�rY��|[�l�����$8(+p��p{�`&�m �V0VKd2HŒ���)�)|��y�m����H�e�:��.+w�Nc��O�*�z���tS�:>߲O�@���3�H�r����E��1��[��E��Ą�`�\OJ4����b�����z�#tq�zP���z�ǭ�)ގ���.�w2�AX.� �k���}m-���C} �d��T�	���6�L��Al����^�M�ocڅ��4������S��q6\:�z*z[>��DN �ٸ��������P�{���p{& �a���@[��<b�`�a֤�$޿X$#���M�[�k$����!�N:� ��2ˋ:�g�=(�B�$yׇ�������ـ ���_���ͳ�$��[��#/��I�@ـ9�*�ͮ��h����Th�!:��n���_��L�O��V�_�8+�+������N�Ȧ�o�G.�j�OŜ�$���Ƒ�Q�Ct砺?%|���)Q�(�*��H�Kխ��")�(�\/R���t����3���.h*�����	�"kKD����FFMx�6�)��hSs��F}G��s��9��%�U���yYMx�ľ��!/ߥ^�ӝ�
���u[�6\݃��X�V�#��wR����\�/�͙���4�k_z�oZ��>���d�q�M-�Z�@M�zH�� �L����X��qe�V��������!��8"�֙�g=�lWZ�.�����.�PwR��E^����Ym�x2�/-��(w7^�p���y�%ǭ2θl��[z�Xy�G�!9�~I��0K6���S�hcM��4dJq��[�p�yg�I3pjȉJ�kMi�*����c�t������BH�ϰW��.�0�m�6�ذ����͇�{H��"�aĹ;{��Pb x�I�����̗((��=})3�ҥ
�7Չ�"DγVY�=՛�B��	Dy���b8�XV�(�����"���2+�T��I�F.�L��d���rq�-=3(<5��L��(L/�"��ѩ�E���qɘ�KG�#��J1��7(���%�'l��ө/��

g�q�]p����&�f̤d��uċ>���,�����m�V�▀~V�����1�5sb��z��m�g�kP��f��<�<�b4����C}�F������r�c=�y|i�S�g�S�|���{���;
֭� �N��ѳX��\,��hr���jR!K �I%k��)�\1��,��v�*�/�.�RfW[��hE,�2�����3�Ho*�ɐa���:-�������Q4&�5�d]����O�E�;`z~��b+�^iE�4����rz�y|�E�1U���q�}�_9t�J�Ȧj�܅��|"`�ћ�C��(�/��b=�N�/�5�}���.��Ԫv2�9Pﻘ��0F
���G<^�e�g�0l�������y���O�,(t���5e�V���[�h���[����2�cXs�5��Y˱��)�H]�by�*�Ź�q���69 U�9����O���2�Xh4�g�D/����A������@ؐ�������j?�������G�p��W�qI�ќXw�?q���í�͞o!t�8H�9�]�[�m�,m��)sC`1�}i�D$�oZf+ӷ�޼���:�(=���c�����3�C��9��1��A��{c7tI�+'l��d�&��ޜ$6��;��x\{M�q����ף\��9JS#}D��i^F9�vM�r~�LN;��	�镻.�a�� �J%T؁a��j8I,k�����I��54��ӆfz�w3u�/���S$�J���D�oC_'ٽ���1΋���J�W��z�_���=5dR�m��z���-C~F��i;�RZ�/�3�`h�R����ohw��4ϤG�=�>�ߣi�<Ne��@r@p�k�����'�La���r�0�/j��1�v�.O1��nm�beă��HwI=�7�4-K�Wϥ��3��M�
�Y��G>����͆\X�(Ց�RO ?�8�tJ�=������ ���O$���^�$z����������}�}Q���_��C�Y�rԤ�FS�l��7^0��Dn�����c?b��?�l������1o�O�
�|UsZUƈ��2E���q�*���܀���hA�Y��&�,r�S@���^/2�e�p2g��;�\��4�"<S����B$&��*��s?^���D=�Ng�2Us@�k�o�,��|��]xn��JY�~|Z�s�g W�뵼��/�g�h?m^�ن�������'e��r!xuQ�]v:-��I���~	ljrU,H�K���"
e2�X��b;B#Qǃ�B�r���
Ф\�͓'�KOk��������?���6�9�)�1��D�?g�ʏ�n�����ۆ����o�qO�j��:�Lƒ�_�v߰t���{6��������˸%~^��{�6�a��F��%[���y��R�F�%�;����H�Q��(�:(��[x�\�)��D;����.���L&F�*������)���^8U�N4� d�����s�|(R!��
U���<�)���8��]p(8<�)�w��(��O��������1�WV(�*�C��%_����(H;773�f\�mq7TE$}Cؒ�����}ܠy�b�2��	{�Jxj��7l# ��7�w;Lu�����Ԛ&y�jN�1�;�ζ�/�]�U:;�� ������C/БT���Fzx��T�f?��؍K!�-������l'ÞW޲�w_��
�n�_���r�B�Y��g����y���U�S���z��5ZG�D���Ji���~�����D`U�Z�w��i���zd�8y]m���*j���x�E�A&ɍȄ;5�r�ys_�9諽�caA�"��eqP��|ǭ=3�2`����`�M��\
�~4Bk�xĈ��>.:�)��dXǄOx��dDf�9x2g��Xl���%�g��qۋrJ�|f|8�(�����/�/�(Ήz/��Bc����x+�+W{�[|�����M�-,Cԧ�G�^V9}9�S�3N�	�	���X��6���Ӿ3��ޖ�'t�����6���a�����S/���[Y@9��~�6�C�q��B&#��#� F��K?�-�K��p#0�ۗ�k���?�krw�txEM�i��]m��	�P���~��7��.����(�^����-�����*���F�o�7l_ȋq�⚦�.^�E� ��c@�5B�������`�u�c�X\vk^��fV�����Eǹ�dY����g>�v��?����+������-A+"	t��׭��/��ߧ��
�ΐA�n;hZ�����XS �rJ(G�T�?�{i�&�Ҹ��_(�8���Y1y?X:�T�.R�lr����-	.��6`͸L�  �j�Kr��>Z>�e�'i$�&��KU����P#њ����������A���H��p�����r�b���_�	Q(�Xz�76�ky�n�	��Z�I[ +vp)�
����e���������P�	%~���Ē�f�6�1�c������]Z6�,R:���r`�o� ϸ�py��n9'�Iv�+�5a����ahHl�]�Dɘ�#7?86�;�p98#�8.}�8���wa��b%���6�Z5rj�z���S rR��6�Є���u�P`�c�f�#����`w�yǔ���=#ɚ�k�[b5a��_v7˞�=t��:�hp�l/	���V_3Nk�y,D��uB�>�Юz�Й�^�0��NR@��7�~��IC �O���
�jqOM�z��j��f�'�#��^�+�6���S4������	��$D#��zP0/���$�2<(31�݌h������Z�c};[��f!����s5`�r8<�
�H�,&��Ӥ��o��t��.�w�Qs�#��]�T?���|Z\��x6B����\�Ϧ+�_���¢�l��e���q�*�����U��v���[mx��Gˆx��m;,��=A��"���V���b��Wr9��ؼ
��&f��E8����2h��G���p)Nk���Ma��|���#�_�>C-��q���L�y^��fm�5��5!����ؤ����W^ݦ��w�,"�`\�T���%��	���^�&��W6�� f�ԈEp=�ȓ�?L�8��g��!�7ED~�(x�Q`�x��G̹���mX��5G1g���M]{�g��J��f���m3��y, Ri���	��8?��$��s��jm��ή�� ��	����E���)u��7+��Ol1��E>=�[^��݊S��a��>f�o�wз�hY�Z!�V�,ky��Uf)偆]�C��q'n��mE��*�0��<kl���a�yY)Td�w��T�n�6������tFC�kkN �>�������q0�m6�Ѱ�4�3���C��XR^�eհ��F-*C�EY��2�	`�g ��T(qńp� ϐ�����5��B[auM��N�>q�W�8��ƿT�t�$�jxy�L�<�*�ۜ���
���[��OŢ��͌���`Bᕞ��� _������(��\n]pK����/.�[�	#��%x�!4��)Cs�����kj�T��ϦȦ�T��RW%bk(VH�5��j�x�2��5^��������a7����FZ����ܒ^���nn��C��?
e�������Hu�h�2��A��Mi�QثG���! �a��j�&گ�e���#�a��e�jjP�G��8<��Ay�+������z���0���@j�j�/������o7W��&沒3a�.���qke�K2�_���"�Dx=�꽢!�Q���O�nS��|�U�ՠg�^4if�T�A����=�Z�_P8:g����!��M{>�:[�~iY�FA؆`�F}����G|�׊�Y��P,��2Vj_
Z;V �j���������AM@�B)�u1��HN��D�+x�"Ξ��(��V���mq�9,���������w����20Ņ\�ҳ��4nb|Ϡ(
0~�2a^��Z�bC��(������4����k�ߧ��3��|ɒ�ZZz��鶺�g���]� ��=C���e� �1[�s���$�<��x����"r���i��҄Ʉ�"9�[Y���a�KN]�C��,0�ubv�_W�Õ��|g�y��؀�2<m�#�$!���jR�tT��f����!(�uJ[��ך~z���F�Eƥ�!��x`�3ׯa��r�eĵ�MCC����ŉ�%���%�e}ڃ���/�s�M������,}�J��*�����[覐<�"��T�'�f���{#��j�����L�)�.C�J^=��U�;������@�K�۽R~�c�,�9

c0n˲k �X�"ԯ�{=�N��ެ�a�`ce������GW�����[/A(�s�"��^: i�{��\nr��o�,�Wn)�?c����������*���	�O���u�,�>\	�2����ބb�7�;,�3�5����%�s`є��k�x��4��Y]����-W!5�Z0JٴLS�w3��\�9�Fa%�LXlxVHYEB    6184     f80�g�@��b��W�Jՙwg��넚F�fv���Ai�`�~0e�Ha+xVZ	M��Þ���t{�lG����@�u����\� �SC��lr�������ADCc�U7.�|�����_q9��^�=ɞN}F�f$�dm�#���>�Sl�uȖ�qD�bޭ>�i�O�W����UBb���YH�7�d4ٸ���{��A���&Y��ZY� 4Q��}��o��y���fv~9A��>c��<iuz�Ao$��t�b���#e#`G&L�<���[��`�)����@��t6�.l�E�X�{��N���"Wr��&Z��d���{�D�!M�,f�D���ٻ6��ſ�e�բi{�5D�J�͔s5��R█����׎d�k;����b���!�;+L2v�E����*�d xԀ�A<:��~�V:�5%,����}�����`�ڤ��9Sx^ γ���+��-��?�= �:/|�5���y� �Q�p��R����M�J�_ X��9����h�K5�]�����3h���O�C��^�VQ�
st��l�]B�$�V��vT-*}�Uċ�+��JC�?�nvu/6��k����!xJPx�i�G�Ͳ�I�
�k儷�z����ݮ���(�� ؗ�<Ϻ���w�i�A��������ρ��k��L�0���l���������K�y��ZS(��]2B|�@I����ȋ����8^�"*�a�RL��Ȋ�}����߃xG�94'�f°�XN9?�.�}�͚��N�A�f���/�f�a�����4�	��FU�L�%<�Tx����W@+L�y1��5�
��*�d�������M���U�LPi�D$�C2�@\`��!�)(�)4�#����%�U�rMT�w�iw�|o���q�YN+)dCt���h@6?iw�;��]m<ٯ�l�Pn��}*
Q�p0���~��+�$u�/��yԶ6���E����Ϣ責6�Ľ�ʵ�c�"V�ڠp�,�cjd�ű���|�sV\Z����7�A�?PA��g$�D:��`�93���ֿq ��E9GSǧ�"	>�6vA���ř��D[�� ���ԅ�� �G��Tl��=�4���1?�<�f�	���T=��-��M}s	�@�.�Q����\jd��A#w���7����-���L����Lp�W �M6�+�Op��aʔD�w��^��3�WAk�yK�� G���.��a��Oe�f���(5r��J�Y��öb8a��Fr����IC!�9���2�xZ�؈�Ue	~7̢�Zp��Y_H�42�H�����qs���cw��[���*u���²�~����ƀ"Ʋ��+�ѫ"8R� =>Bk�ӫ��c�N>����=~A{Q{�fs�Z>_�C�ə�N����\�-cc���pG�	o�hx�q�1�Î��r�q� ..zR��v�� sx)���AxA+:�MSg,�3�v������U��=M j;f��Y%M�e	 �a2.{s�'Zc&[4nw�SLQ�ܛJ ۦȁ��If��m1�������(��KmB�����כ��^ܧ�*�~��q铽m�ǅ|�w�t�������U�7~���ص�h�g��"e2:� ���H���2:�฼�Blʣ�W�����:@Q>n��= J�,g�3�f[}����6�p�m�;m|ytx����8��p�]Ҋ�]�[���q]�������T�	���B,�,-���_4U$�v�@���el��93w�)T��U�6���2S�a6%� ���3���IK�O��P[���39Q��Z+ �yF������`�G���`t�4�V��^ܯ[?��bwf��w[t���]24���{�2����nc�2z��
�čy��թ�s�crr:�'܈���kU5$�t��"6a���}Q!;a=ceqUv�B	�eXߡ�;���s`g^\+�b�1Um�"60�����9���qb6�E[/��O�EϠ��A���X-h�������u	?�!e�����o��0@����h;GXh��ת_{�h������p�r�^��0��'.r���.y&�j�]�/�Z��?�pʫ���]y��r�Lw&΢#6�Y�1?���̓��)>�h#���N�y]c&��5�cSj�▉'_��$�����r|��f���78׽�&(�y�*n��	�4W?<�z�HE�	�/_�ƽ�~J��tP�V>�=�x��TE�$�� ���*N� MlA#	%�Ѡ�,�I i�a��Y;=ѿ����ůM;�18v��XH���
la�2�����%Z��\�d��E�݃������]�+��[�ė���bj�<��DG9��c)�n���=�(�a�x2�g�\�z
Z`x��(6N�dN���mTwǏ<��V�j��N�d�MO���2q�n*�i��-[�J���7�|�R�R+w#}<��E���DPVyu��/�hstYۛ����ɉ��́2�D�S���}����hFݽ�&-���h��+~T��>��sAb^�<+���Dnp �4��2B\L�^B-���25\��Di���z�3
�8�9\G��|���	u[��,�g-�Ơ|D�9qR�k�7f;p`3��_1L���bN�
�9{�J�֛���ׂ��� ^B~گ�)�WƎ��M����]W��@�`�$�s��@�/C��y��h�����%/7�{˕�hSs�(���t�@��BC�dʈ�Mpc�<p�*ױJ���(�1��5�`:V?�@��q���K++rp�p/Thu�8;�,Mk�:E8S[��Ԧ��j��$+�n�9D�G�a:0� 5��c��$�0�3��'(1|ɾ��; ~��N����R��5�����?�Z�I��n'�ҷ��os�4��V�un/$P�"����*/�;��G����x�~�.$EHG4W<�I����1�;���Ya ?����x���oߟ��3x�E�W�{�3�3V~�����낺����=�@r� �����1� . j$�E�P)����r��	p{f;�+ �"�U�PG���в��s#�.��@�ů��CW�̿�w�d�3Y�35���[l�I	�Vx�&�����d����C�m�~0_�h>����{�}{x�Й8��g[�-�o8��m�V���;��������b�}a�����Y�r�}Y�n��H��q�D��Y��T��oă�h����Y� %�/�?�|#�o�C'��bq�mеysuL
��<�8��jEHi����=
����V\9��6V���f�4U�-���l���2_��u?��o*�]���$�	[�Wȟ��z�瘢T0�P3@�ꑳ�DX���x��v�*
|3*Y=&�:c2'15}G�����s��*|�$1�G�Km��A0��D�����*��/R2{�k9d�Z�pP����k����2�8r��FS	%� 1���xb����aɲhK��if^�V�F�{u����d�^⩁���M�?�����˽�A 2�d�'�������`�<��O�i�l�4���?e��&ɘ�-oRV3��[�j@Hp���'y*D5���k	4Ͱ��fZ�䧣Ed��s7T����xԠ%�NA(��~�A���/sM��'F�M����[I�x=�Ŗ��h
�O���T��+5}�"����D�oô��I�&��r����%*�Fl�'N��M\Y`��j��a�LI�윽�a�uU1<^��G׆5���Z\>􉇮j�J�'�9�֦�G�_҂�7���,@o`�9�u��M��
]����8��Kה��0,[������=�Eυj�Oy���n19�����o��Ht����6�_屃��W�Wm��h���:��y�HÝRMO&�=�t���{џq1*ռ���j'/� �f_|{ 