XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���haE��GTi[�{C�;ėU�K�B_A������n[�հ�FЄ�3�!��),#��[�M�/J���<v���d ���Vf4��������bߛ3�JR�zC9�d���q8;ð(Ae�T�T1̿�͗H}�����y��9�Emp&?x�(Gk9���t\��c3<P���!2�����u.)A���I#>���O���l=�_p�15}if,��)ɕ����@}��O�-��I&���*q�ƹ�����г�'	��TW�'HZ�"`��8��t }[h[?�����L���ƥ�������B���E�T�m�8�H�S ux�~���(�-|
 �H6-�����F<Y������C��U[�����}���@��H9I��n��о��'����(���hMP-	5������glt
hOn޻�]�rNP�X�����7T���I�n�N� �x�3��dyYg�M�.�H.;��t�����^�����#��G�H�i�u�q~��R�2r�|��*	o�Gֲ��C	���0�R,\���Bؙ���y�+�lj���=<0��Iq���X�id4���U2¦Z����l����V�N�A�?� �6�6�*�ex�p(���'&]�v_��ܷ���,���0(���=�X���VUR?o����H�fP<�~r1g^�����3O_�w]-��R�u�|���d|n�П��I���,�1�VXch�^�Ң��dKi����s�z�.��XlxVHYEB    162c     850m/	���Rd�QԬG=9�7�L�"E��ԫ1�Nu��9v-m��3R#Gnڴ7�����d��B��i�;NR{Pۖ��y�LL|H6�/�M�%�@��f��U�tHo#t[��]n���M�Ó�]xU��ӳ��Sh����&���U����X|5ٹ��`�W�"��Zr��O��ht|�kء�mu�F"��,����(i\��{��a�`���;9�Q{N���(��]�^����߭�mG��.��ܞ���<a����!Yl1�p��uU;d��@\G߳WF�L��꾡�*Fqy5-���ʘS]:�?/�zY!������ƭ0�P!
rJYj��F]|DW���͡�j��T�O-̮E{R�y�0vöo�@LKۍ/��5I�}@��d����Q[!�tkbb�?qƂ�z���۷�}�rȭ���׺\�ׇ�J�i",��!|�H����_0��&�8�����5?����sz�YM�k���d����7\�fˀ��w�+��q�`!�I�/E��sQ��&'��Zxߑ��Cw�x�~����a���gO Ա�/��]��7$��W�����ƆT3�D�fX��Y�@����e���᳒ן�#1PcP�-YU{7 i����lVhe?H@����~�dW�H���D�[�"O#����W�,h7��V�6�Ni��9�X������8|�w��^6�#��[���E���<�*�m<��⼸X�ݼ���t��νIa�*7$�+����͑��j3��tlM�,��_��<	�mW�Gm��`Y���a�x��ߴp��'��o)�~`�d��{�B��0�si%x#QM�y��U饁���#�`��>C�T}�*������f%��/�H,f`���䌡Z��9���u����1�����(�DQZHi`�@9~�ՙb%�cEڳT�l���E���dG�'v&¤�s�c��� :!������C���G��K�.]	�mY��Le����p�w5�7�d��I��н�����yɨ�%��V&��v⥳9�DV,Ӝ�o>�8XaT0�֬v6	�}鎜������"������<�����ͼ����9��It+�e��h����(����c��H��t��K��,�.�MB_����J4��ѦC�>#9�Rk�΃�#�����K���ϧ`��=���zT>L�5��5s��O��L�\��횔������}R������Ǽ����G~l���P
"'n�)�	�s"H.�+����Bω��3^���p��+D�:圀 �[Q���t1z�Wvp�HnO�|'����`3Ri}�_��zՠֳ���S���)�E0̈d���,��8��&P	���:�4�T|~��
��T��S[�+�.8^�bQg�Ⱥ��%do�6	�̈́,C�PC��Ks,�r�-���#�i�'����W���]���L�b8V����d���C���ᅂ5%���݂��oު@�+�|�<g����S���f��b�AGo9��~�&,2�u�@�C��ak\Bո����Q=��"�)>��C)�2���^�l>a%t���J���2:V(����'L�<U�7S��-:�"|��v�Y@�tX?i�j�����N�y�����nd�y��W�����Y�^D��9�Q�� �zWiE�i��^�؊������ͅƲA��)0���q�PqX�������;�D�]����e7�zְsWހ�E��,ekqL��f ��[��|��2�C6�ś�rR𿵟X~�l�XN��S�Q-���@5U���� '���P��\mG*���K����ȟ������"�6�K����
��	�<ƣa���%��i���En��mA��i���Aa3x6n�ۃ}�b��qд���0�I��@��b��,"��O���Տ÷|����q�C��uٌ��o��;��Hi����g&�����lz�f��򷼽:��L�	��=lڥZ�}�, �ע~G�@߾��	v_?�V�i�n�/9T�H�6�en�`�ñäػA��.���8Q.IU��p#��7��,��y쑶m8�2(��gU���