XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%��7B�f�D�֦9b`{<�E��Z�Q$����CO��_�jY@�Q�S7����i>A�{47�1�}$����^ǽ��Ti�A8loE�&��d~x|����5xu����
# �Q�<��N%|sEh~�a*Gx��w��1}����C{q�'�:{z'I`p�6p�n�ݱʵo����F�d�sZ�2&Vk(x�|r�I��k�k���t��n�,->v��9{q���]B`9qiݱh"�>
e�5>x�m��L*������rJo�dZ"�;��[�`�j����v�"�����+%|e+�j:Q�ߪ�vg�CR��t-�L�֧=��թ���Ba�O֓Ԗ�m6�KV�1=QduH�	%P�1ǌ��7��>���f���Ir�2ߕ>,02?�y%��i����$)9+N~�����^�Ŵ���S�g�hQ�-��7�B{�ku���b���m��T��HW�nM�z��ם BI�˯�6{�[�]oЎʾ�m=ԟ)��;Por	��-�޻�!�w)�(`�M}6d��0�)���X�Kk�>0>#y[�O����~]%��ӌ�|��p׋�U�=$�n�#��<��2���4��2���� qyp[6�[W�(�
s���z�r���U�4G����'�'SL`:�@���Q���l�Z��b}>��4"Ӊ���WoȨ]��?9��*@���K�$�/}��Ɠ�Ͱ�p���{��M�̠�ܞD
�c�0Wڟx��K��bgL
ËXlxVHYEB    fa00    2950�,7+Ez�ߥO@g;ɼ5�X�(�c��W��ⷔ�������y�[(�(p�,�I��䂏Χ]��p�m���L�������Dw���F �e��0���3e��c3 ^cQ@��cf��������T�|�=mtL�W�1c��V�̶�v�W�?�k�Å� �Y��~�.�G�ر�7_U��Ȑ\N�¬�FY�]�E+�`S$F:uݱwas�W��U�D�I��sG�(�õ�e�82�9� �5�Bo����Q��}b��B�h�%�ch����4��`���m�*q!���Dr�as~۱
a��>�)��?�?8zl�:˛;혽�L��Gds�����6*��]��fҴ��R8�݈\y���F���d>lse�}D�C#��(������W��^���E���:�m��a�8��89S��?�5���k�����r��\��N��h�։�jI�c�
�	�Y�'*<���t3~�45�_�:�	��Nk�I��`����%d%��!�R��>�y�{��)�_Ժ)�z��K�����|j֙&�Gܱ�׀d�BS@��G��oa�)%̙}�u`��@vz�X��'�����?�)|- �?�5�.O�����K1cpu�=S[��i�=�~��k�4.W>�r�:�Q%�i&~�	�1�!\�9�5a7Ϩ�Y�Ԅ@�/>��k9��'��<jg�a�)sj#X\���p���]'f��� ��CP�zˊ����'H�gu���MA<�Ҝ"��e�Uo�1�,��䏳��h��T{N������R���?���\ɴ�g��aJ�K��A�"	k���J׌���E��uݯ[U_��	�����/�I��>���Ցy���"�b
���$Q�s��4��<}�����$\��ˊ�O���'.E#4C�I�w����5����;"������V�d�娿�/�����������~����!�~�q�YĤ4��iߢ�]$ �y����/O��D.?S �jY珼��Pf;�A&|���*�m�k��]z��c1�����o�3��Ҵ'C�0�iғ���˲]o�U�I�v,��Y���>����5�z���a��D�L��S�
2�(����[��̳|�����`B��]o���A4em4NTV�P������%0���74�|$��E'$L���}�}Gp����Gn��k��R��Co�S��}G�'�?���ϼw��jyC�b9<<��Pʛg-�AZ�Rn�M9и���Zٸ���Dȵ�,�9�Y��H <�~qh����oy�w
IJ����-��Y�}�2�:�����ΕS�V�%�1�qs�O=>�?���U�E>H���P(
oQ���xP�Q�K`	���t��42z�"���	o�	p|�#�Ā�25��i����hC�m?Y�&���G}��+�-R�Y^	w6S�Dڷ;Ų�56VB_L�3�^������7�t��N�9���eL]+��Yr_�(�����Rp@
}��'F M�Fn
5�`s�b6����+v�C3B͖�8��#�=�p<JU�%����C�x��D� ���G�H\QV$��~ ����ß;�G� ����#D�\<��@�������a���`������u� ��|�g�l�'VO�BLO
����\��ː@�V3l"x�-(� D�_��A���TD�#b�{ �����1�ݐJ}�+�SqKQ�\�?ƛ�
���� ������̎��k����L����m����z�Z��k�+�+���.$�@�4���ԁ�o�c�Y JN������3���^�����1�p�D�"C��� ��X��6���0	�0��0PG��2 ��G+�%ޒ�N�g���~%��0�9�
U�37(�e^.E�XA�cj�R�"����:Tvyf�G�����y��4|ׄn���������$s$*QR��Mh)UwX�>�#����W���c���\ɿ+�m��C��*Ǉ�.�ؘ}��b�Iw�J'k.S��Co�$���cGc&�CԞ��kq��c�@[�k������}�uQ-\���
���9os���''Sd��mb�=s�!�i�?�����gO]I�p�B�������������w���{��Գ��.�N���tJK\���K�'*�U������ͫ�f��>E������ �[5Y{��W��������]Z��e�H=	�kVZE�l��Ak����4C`r74�s���_��o�a���Z��Ƞ��6�h9�?<S�
%g��H�z�}���<�HąG �{n�*��V��d��\��k���,ϟ\�Hgu+ҽ��d��l�;�&ϲ������N���&s <��r����TG=�z0E�e3�����gA�~�^J�A�o��B-9k�\��o�-��� l=��E�*%�2t��K�Y� �}�]��L]Tx����GD��$�)�,W�$��!���KOlV���p#8�˅���s�F	��}X��h�g�$ŮR�1M���'V���|���d犈bh��)nW�E$��d1`�u�c7�9���PpA�VIĄU�Ť�K_��:�ֿ?�9�)4�||�Y�~-��e�0o �/���,b������f4�a��Wc�ڿ6H����2 J��<Y<e:��CVd>|1t�R�cMH�a�'�A��-���D*�g��� Im�r���?ߺ��LAh@u��Z�ʜ���C-L���+��OE=/|��o.����
R���]܁�IvE*�tܶ yE��f��o >o�q�U�����Z�o�N�ֺ�C;<�Xc�`�9޼7�	�wΜw���%�}�[�u��z)�As����.;IA�-"�}�f�7��"�M�2��p�Qn��U�k\���j�	[�o��A��I�>$�r�-�p��σ��/��_;�/�͘,��Dc[�k[MH�t�'5�+�����̶1�ɩ.3�ڿ�щN�2\*��f��/�u���$��8�04X�SgQqZ����A{\����Z�z�[��[���lt�.�!�垈L:SQz�%O�5H�׋���u5����|����(�G?����"����昆�ե�p2�4����i����6����@�>���@&|v�C���N���V:�as?Jc��B2��dd�G�j�������O�UN�9�::3i+HY;�R�3�-T��-����!���:+H��-�)�R�n�F킈���q�� }�J����
9���u ���̎���N_��,7��6̀.8?�N�
��5���NhQ/�����? :�o�[^�?�G��`�[���4c$�ȝi
����c��དS��=^�L�ն��&d.����׻�+��ՠB�Pnu���.�L�N��z�*xL����M'���6!��#p��;j�Ȃ2d�=�B�d���z�R�]|�@'�#����o+v�`�}3l�F�%��bomn�!r�.��G��'���颓B�9�� ��qh:�=��XL�G����7��Qԫ��N��y�N?�˚�'��pV��m�q8eL�	��u���˺p��ph��l��Xk�9������5��a���xO���u��V_zz2G<����2$��t)��0�8&�H�3p8�l��Ym�j�D�t��֧����=7=gP�)�FD��Z�G"�G�K骢�)<(uB4�3F	��巽�b���)�`��H��m�l�ҽ��+�?�b��:��Y`�ʅ�������{cl�a�0�O�]XB�],��p�;R�WA�Pvu��lE�OÄ`7[�Ha���"��c�n����f �6�QyC:�yfD��gg*��8a��ߖL�L|m^/�=%��*驧<B�����u_[����8Gf��}k�up���]}�@�z:���)ϑ1h����s�/N�0|NA�넻i
6^�X��]G�5|���"v�,�����2ʍ��\Sa��^=r��N�q��`	 ��2d�����_�W��3a*[�1���>y����IS���.A�����ʾF]0I�|����+W!�J�V�F:���_uJ1�?8F��i��/Uv�&�[�m�2�nI�P�|�>b�v��{���ʋ(�,KV��$0����>�	�����`` 0Ι/c\bJe�>�g�K�����(��?W���}y&��E�	m�"zب�O��0)z #���Pj-*�:��Z)�KB�n�eM|&� ̼�����;K`q]z
���,g�^*����/m��A���E D4�6��og2qK�n�Z��x��J�z���O@Y�?�Ԏ��ؿ��W���i:�3�3 �}�<�=h4J�G/�'IN�1��/(Fa�~�I��8*j_r�S����-�M��`?�����ƻ��jKg�=�	,uA��S�g��=�JJ"��oL��D��5o]�'d�P�t����pg�Z9z�xl��Q�#ז�;.4\�>��g�zy�En����N4�4tF蕲�6�v��Jv�,�B�O@��*t�қ�jC� P�敌]���P�@j5Z��=���*6U4 �h�j�.1}��nX�>�@� O�����_G�֚�:ǝ��Wo�<�p���Q�^����Q�O�qg���~�'�\��8��-��#a����L��h%m�Js��'�gi�����x��>���\1�IR�ۯӲ�X1����U�&�y��W-�仯��83�ՋNw~�= ��!l���/D'#>�S����e!��:Ka�(K�(]#�%e�ԭ7E�z#h
��?Ic�(pmE|:��C��ւL╅�ڢ��T��Zz������6_�������OX.����H�����t�ˏ�\�h��R��(�Uz?��3�!���q����8�5��?�	���	x�1��Sr�-_p�} uh��7�I<�wPx��i��P���B�����N���a/l����w:/)��a7����I�?�)d�iެ�e�w��o�%�Q ǐs,�^�}߲N�~�1-e)��o������<���� �o�f�UP�9�,RT)y#
_�+`��gpz���*W�e�W�[���֥��-ԉ��N�����!E�0���[�pE@^�ƴ]#?�յ�!/� �翟�'�%�@
�G�e�.��Ĳ/��ݼ���x�X�>��^��hP/��j́��#�F\�࠷�on;K�g��Μ݊f$K9�
x��̳� *�+<���(�9��/_�!O=)�goW���I��)�վ�v��t�_�Э�!�	�ʝV�d'�0�uc$"Uݩc%@�P�𬂭�;܉��3{��7�b2��@!��R3G�%�x��Z��/��ҸO����Ys����`��U�j�����߷O�o�T9�����eg�1-�1��E��[_��T�C��V��������������o��ڿxR#O�.-˖1�Z
�[�a$�4]Y����(����h�M1.���a��;Hr�E}�b��� 7|T�&\����bK�떭�P�m���B`����r/���gc��Cu�fD����ϯl߿��Mr�s�$]H���XМA
/�ػ=>��VX�I��C'XL֙u`�~��xc�F��M���Z�]�>����n/��4���~z����s��y�����~�P]#��ے�u�ͨWjdZ�i9o����:� $F�C��J�;�mG(�}��`J_hX��3�Bş���;?��VDC���I��ᐖ�[��(C�z�V��5	��d&�r&v�.�w�g��z�)�C��f ǳ�5w	s6@�5����ne�YLW4d�|~��VA�V�۔�B����;�^�h���s-3��hҪ?v������jeF�\. ܀�b���f+W+!�VY7sB�f��J�wL�.#�D��	J���N� ntq$d�E#����Y"��dz"o �[)g�b�����[W��t�a�?62,�cyΕ�B.�GYUiL��a��܀�Ws<����z��6�v�k�d��K�k�U���� R�Ł6B�n�,ٍ&�>���X}k��+�\��Ѝ~�R��������6��yh:D,���U~�X���T�Lr�R?W�E`�s_� ��߈�!�U��On�6���V�p ����e��=�q�rų�n'e�{{�;����1�J�M�wuvb?�f���W�����i���7?�t^�Ye��L��a��d��<�G����U*s�/�2��_y�#<ʒ"��j�K������@V�`����b/q٥��$�;�"�EH��By�@����@%r�E��؃8͗��l3���c��g�
m�|��`\���=��_f�Y.�}���P�Cqp&̒�8�>=+�;;�~,�<��îG����.��6Ǟ�/�@~��
2�hhJ���l!n@vg�M��C�7�K�Ŝ�m��?�**��G��F�ɔ����h ۍ��b*X!�OQO�װA�N����&�n.��g(�
qS���i%{�i��D�����2�K�荷e�2~8������"���}�AC��\iG3r�7bf��97��(7�b⁶�m,Ǳ\j��M¤Res��9�t-��t��<���G�W/@�¢���<n<�B�m(=��CC�]]�$��)�΋7��M��w�7I�W%2W����no96��=)�Ǆ:��Sq	����i��2}z�R��ER����S��ك�V��Hɯ� ��x��a>+B���o�pM����jT%I&�Ћ'yE������f[���-��yO��@�>Wםm�x�(��ۃ��l���l���O���L�� �@u����@rw>/ �hk��������U�uc�?�c���)S5AZ�T[	%��IP�"��W~i���i�&��y�b]f�t�������+?
5ѽ7��Sp����݂�;�&����s{j�� �~�T�A/�勀���`�����+c�����ї�1�ʱ�H
�i����r2&s��M�`�`�0΂�6�O���9-dˈ���7j`O���V��	/F��/�8�E��|y`�SF��t|�B� -���sDJ�׍~����$�z��0��lv	blB���RWg�]��i�ɉ�9�5m���� K�ݑD��UL��&��:�J��N��Y�~���7�� ���q�K/I�mA1{Y$�C] 埚MN���'j�t	@Ǐ�n0�"I�V�)7=yǪ�������)��bA�������{@�w��դi�Y\�>8��eZ�o�rAa��Õ�-Rڠ���5f��9@A��ڹ��v������%��&(A���o�	��Ua�����8�QZ^�w䫪��N����B����o;���1�n�o��f��ة�>�I0h�` ��@�Wk�Yn<o��c�����]�rV��#����~	�Ϯ�=}|��S2�F�'s���逶���a��$Tf��������KX*?p4����쟦�f���31c]{e%���e_�Y��5�L��;�4lT���B�ъ}�e�?%1��������q�'x�T�Hg�~7���`�ꔄ����/�Ox�����[�R�0#�c�ky���=ܲ�;�R?�t����=�wU�;�Q!SW�t�ǌ$喨j�����-�R5 ��X]����	�K�E/?oA��N�~W
����N"���TsAa���%�;�F�G��$��c�{�Wi_���=2���ۼp��q	� ):�����D-����G�DP�K��V��$;ɵ�f��O
rt8"13�o�}�xL��]��8c��.J��U`���f�܀VW��5Ί�#��2�+�ؘ���9$v6}���Ô�έG@>t{�cub�x�%켭ws��P� �qq��u�v�5x��/���U	U�[�P�[=���EaR���E�^��Ah����3S���mϤg�趬]�;g4���_��_���K��o}=�vcyJs^�K�'���s���	��.�̈�Ub��9*�2��b�陭��]ٽͬI\-	�B�AJ�	�"��	v��H�mqIs�6A�?�Q8�]�/�]�Mbu��l�qs���<�T(���ށy�vW�B��Y�vM=@�� �V
���C343-�J�4�tHJ��p��W�����B	z��)�U�*ƙ�J~S���W��-#u�eg&����D�-����"�Y���y�V�|�J��9\�Am��<t��u�_��!lr �x���.bv,F!�*�! ?b����ۅFL�.�Κ�>�4��)p���)\��D�~,zL���>�q��On��m�:�vmAp���g��_ �?���-�������)���@$�ka
f.��Sű+S^^������Q�	�_��+�*܆�;c\O�L��n9���.Q(Z��!zi���Eڸ�aIM�ϐ������c�}�� �dL���Kњ%&���E	���'2�?ׯ$w���$��2on� �KҔ����*߾Ѳ�W�5Ϝ���v��Ƈ�y�^� �~�uq����c�i�M�'⽊/�WI܆�l,j���8������=�⍃��!!cIڅZO�9,���M��u��7f9r��߲t��W�gD��Y��T��%zIP�d�3�"k�(�����yA< �/9��lo��a�(CT�V@���Oq�,w�m�[���	�:�����Y����2��A�#k�#�#�e�կ�Ir��H��D���Y	nWVmҐV1��z������x-�BfM���|��=R1X�Rӕ����p��adzN*S+sAi��:�>�����Q���솱@ϱH:tn�� �(�1WY:��V��;NX��dZ�}3� ��6�zA���j�«��y"�C�E�b��<J������d�J�PJ��ô�"$|���7;O�B��_�zP�}%��^1�#	:y��͉�}��Z#L�K�p�T�� ���rj�����AbxU�)6*w6B��-ZfF7j��	�u'�u�}���#���13|�ȹB�) 0�(��[nkxy��+���e���$3ɸ�#�q:)87��&j��J98Y��xX3��
]����'*
V7ZΟiv�W�����F�tq>�rH���6L�=�M�b	P𶷒�n��up��2��&ֽb�Խ���V_�%̬�r4�:S�����(?C�]�&w�������GKu>���U�r����x�9��= =��(���%T��p�:�fc�Ē��L������tlR/<j�	F(��/�g8�]�Y�����dEi�H���a�`M�/-��+��o�s=G)��QA�5n!m�e�
��*�<I<9���(A�UbW��V�ᯪn��ƻ�����5W��$��/��,��S�[�;�#�^����0�}A(�v!>���t��ܞ��0�W*���*��E@�hh�� ����W#9^w`f�� $��<8�[���:��� �1x�E��֫���?�<l��#�v^l�vr�����_���_���I�+i
o_C��E9	���5�,��������o���9�D��;U��l�����L�Βޜ�C��j/�&6;�Q�t���1��JP{��+�(���ԼmM���H,����,#O��dk.V=k�}��'�wa�,ޡeaUEL�\�ԓ�@����Xܳ�
�"h?L D&ŨL��8� �U���Hɑ-݋?2�QE˩x��Y����d�/�U�Dco�_�JR.�5kr�(��2���"%"���Z�ߥ�;��|��Ng�"ɟ���*�z#�?��g�e)�Y�:@k�8�
��O����sM�~��ތ!v�S��KN��q=[�̙c�E��bao\��?j��׹�أ�i�9�����Pu�hG�0'��hp�����,Ӌ�{:��)X��D�<T27%���'����	�:{���L� ����ySĥ����0_I2����ZW`b��M�����_r8grhD�)�Y��~u�=���X������*�Ǡ`�&�&kx�ܟ��\B ��~`������hn�},�R15����p�aN����>o���u���̨F�kG�Y���+��׹uz�B�����MZ\�;� ��7�`F�8��C�{��o��T��a����^g��L�_ϐfH+����h4��m���e� mrW�o��ťїxEE>X�V+�����ٙ�*q�,U�oU��Qdg�i��V�h�����_+�{�݉�8���G@����Ș�`�|��[�#�����i� ����0H��f:����f��ae���^�q��a�B32֏
w�U�
�H'��w�bQ��	L�՚�L��ecUD]�>-_`xx;3B�w��z� ��(���r~#cD����mK�#=XlxVHYEB    fa00    1e30+م�����<*��m�A�����c�$�|�*�"�n_�ߊ6��G�`���&���i�)˶�����c��a@�����(���&��|�d��:���d�2��R)_�2���W��?��ǖ叓�
S�I�����fc�����^�j��1��T�k�9�`m�pj
�r����ߛ��0ȢT�1��'��OƑC��ģ_Fږb���x�tc��KCڜ@�_T���W�1%^y���y�ζ/Rn%5E� u�^�K��&�Nl����}�.�2-u��iG�<��������<�YA+�$��A��������#`y&����n��c���#�wyW���G�s87^~E&�t#xu�p�ͺ#퉤;N�PW��$8����R�5\�Cȟ������N�WyW���1�hE�"��	�@�����HD���t�q79���#8&�tA��21cͼ-�L}�\\�ը{��G')�f�g���!�l*b>�n�i5��vuIn��	��X˱aa\���^��	��w�=�bI��&�_*k��\����� (f���=?_��=����$"rXf7�J.�_���Ü�:Ov�S|t��O^ߙb��,RݹUs��Bƽ���?>���b�N��:f^����'0xGۓ_fqa'�L��o�h��δ)CB>Fn����9)�����mKM�!I}_�4����Y��u� ޱR�rK�°��"bP�[��ށ1L��9 �!i\��}8";t�ƲI���H�Ӗ�k��zn䚶]� Ƥrmbw�R ��F�׼�#��h!����7D�&�:s��9&6+�1X{ج��%~��AX��b,�	��gh�9�.�̋�ed�bbb�%9FcG�!%L��/I�?�dM� ױЇ�<��|�{'�cG$fe����r@×�s���D�/��z����	~�p�Ww<h�`���#'�ܯ�Vg��y	]�{r2	a��Bv�ub^��D d��Lk�K�}����Gr,�-1ל��D4��/c�͝�Dc��)�	�(�9�>!����^=	�̨�}Y��3�x�4�x"�b쿻+�r�����;Χ�6�v�J!��^������fb� "D�l	�OWCD܇����P��0s��1������:��c<bE3N��en�X\�c��Mq��H�":KQe���p�l�
���u���T	��*[#dr�ǒ	h�|�8rZ:Cm����H�g�;��MŽ�dR���~fU���z��n^d/��W~'�X�1�F0�(�4����������H�X�%��:%�I�C�fB�d�m�p�����-��~3e��2)!$;�?oq�m�E�(�F����dmAy���|=�������ы@<'�X�>�	kK���~仱����P�"<1E�޾iyhX����9?ӻb�ۉ�(�l�����߀W�){�d� �eG�\��V9M��U���aϺ��䚚�lD���ÞPG{dq�|%�c�J��-��ĭ����/t�!��-2.N�<��BJ�\����>� Jq��-�g��~�w�N&�=�A��i`��ҟO�^�5��`*���D�����*����ʝ����qz.;oR��=��޸ɵ�ͼ��?����1y�4����-�V��^���j�.↶��p�N ����( d{�Sm|uuԴ�5� ����G�5�Ϲ�=���^���3�j�Fu7L�Hj�w���L�Q��	3����7�)|"K�esm�Z����q�w��!��A#�BF^S�enO�����1��B����$5k@����؎��f�	3�$k�|�����_�2;5u^����v��1J-5ꅋ�b��\�8��	(ߑ�#Ŀ�wƮp@�D�3Ϧ�����R�X��[#�� ������[��7�����֒}x�yk����z"r0�$��+^�+"��͕Ū�|߸�{���A���Y)�a�6�Sg�.�N��8d=���&{��9XqW��Wuv@[)*�R_ϋ%�l�
��ccBp���b`@�h�K�#
�5�l��r܉-]��x5r�b1�HV����s���|&��i�ªtۖ�P����K�U�v��^�� ��������jt�1�u�M^1$��U�r|�͵=��7y�+[��\��/���;�RfU���Z�׺�����F����
�Տ��H�VF�ܕ$��N��	d�n���Q�*,a����Bˁ	|�=��&���'|��AC�*_:U��"K�'J:,�C��V��(�U���v�Eϡ���Kg�!�O�1ƏCaW�pz�'�?���J�ڱ%b\��c���=�%:�:�=����Q���7m8a V�΅<����+�.R��|"
��S����VT"�q��m ﹿ����8]c�Q��쎺Dj�Ԗ3�"$�b�*V3nӼK�槫����0�/��W���ֆ��MP������_=!xeEm5�L"!�������R8��+�]�}�s�C�/�.�	4d9e��y�E�C��{F[����;n�k���ֵ�d����M������2�ԝJ�$[��t4/F�5;�=r���#�1a6c�qñr1� ���<���iO��������o�&E�| �0/����A��R,Fg����l�[Ka(�⢰
��)b,6w�9��)�M�����s�.�f��ύ����Xv[�O�gLo������W�B�y� mGe�C|B�'qG���UE5�ȅ���|m6�e�D�%S�,k���0�����X�,VS�cKoI�=N����7��=}|�W�k��W���7��q��y~��wA��6OR��peـp"J�ʊ��3�@��zʃ�N���S3�Ҕ��P�ڲ7@���� ccr�u�#�-{P511�n*2���#ᄌ"�;ʖ�Wd�\��Kx!`~�OV��z{Z7PC���(���b,;͚�!r#'��`�:��;V�Y��y�^�z��ٸ.���HW��e�=�\u��e\� +@�#�pC���*j8�{$�aԥ�zW�3�%G���Z�.h�e����/Mk�3���?񥐆��}S�4�H+�G�	�jǌ��@oam��5�0�]�4@���E$��@B>��ďŁ:[5G2��<;s�#¥ѿ�e���^�6�n�e��Y�^�m8� �}܈�u7.�!پ>����-$}Cca5:�<w�[�N�I��e�]�'Qߝ���h���w��H&��sm�~|��K(��-^��l/���n*$wl���}õb��x ����O3��S�:�p&p��E-����eת72��S!��'�.j�s��*a��<��u��Q����T_�s���v7�K=���AnK2�:�0�*&��k��l�S�"�-�<X��<z�-x!�VEZ �D�|̏gXc
+�I'���"<e5N�!r9[��qN�a|����n���/���VG���8)Y��5:�s	�ՐͅS"EX���l���_4��;�
�����<t�,����+��^&��bx`���pFȗ��#�<Mm��0��Դrއ6��1k^jWX�qZ�z�`W�zݞ�2��׭Cx��sz�Z�.�]B�̆2O�?�k��]yf�c���-
�aͬ[]p��i��J�ʭː97��N﵂lXb�vzr� NKV4��,�\k��!���#m��n��Сff���:f~�	�~^�0�I�p���9
"����pY��ACM�~���T�_��h�%�U���{mDІ�rD.�9�~a��H�L�o{my��'o���h�a�b����$�Iԍ{��L�k�B&4�XJ�{C/΂��C<.Q�­̹�E3�z�OۣG	�<��
�N��f,V��z�hQj��龷�S��� �I����o�^�=B�^�W%Z23���������s�%�+#1��[�O�NaBԮ833/���j�	>�ƅz[|��A�T?j	��<����u6�jmsK`ש^�������l]�я�:\�K�jr4�4���$��퇍��s
O>������Q��rQl��׬�%�fW24$%�Ո�@���݆��g���@)��n��Ey
(�jgev��(w�1��uQ5� ,K�+|�����j�z���Cjl�Ҏk��a�pзz2%�*0\���l�"���-L�d#�"j?����L����^|nH|a����߀�%x��Z�+?}�Z��{�f�+`?�u}ɐ�2���[�H]4f9�<�_�R��� ��ȭ�m*���פ }KaP[o�v�).M�����ڭ�Ր��~��=����:�L"��1U�/�?H�P��ɑ�Fo!r��e��L$�;�9��5�N�����6�k�m�A��S5��8jCqRoM�rgq�W�����铇o@�,��ukn�ˠ�
�d���C%��kor?���vE����zQ��e�ۘ�U�>Y�M���P)Ծ������@w�B�'R.��)���&�hx���Sa7��w�̳!�I����!�B����)r#*��C��2o���j�7@I8U�"�,9d��c�K~>(�sն�ȇ�*y�E 4{��Ry�ƕ0b�T����d�ӎw�}��-p��X��ҔMp��.�y��)�� ��4��cY��0ck�&x�Z�gw�$X2�h�����<�(���ҩ��PkO)6}L1F-����.�m��4�;!p"|p)�����4~���k�����4� Uk��򩎈�[|�>�����͙�*�����9���1W�I-yHB���& ah|��p�C��V�f���|�,�|�{%+��0�(��d68d� �'����yH0�\��vĨ&�2�%\�{<s6��+�5T��Dv^�ȁ�7��Q�������X(��2��2�\��Si�h���sN�i�{?�B`>�:���ج����- ���Y�u0���Y:ys����=7lƍ|��(���.�<�6:yX�|��Yr
�2� ~V��i�K��D�fV���L�Cn[����t���B8}u�XK%=��r��o`x�5��A�qkV�qB��ە
c�(^�>����<���e�^�P���4!��\�+�T�Z��-����V]�nc�6@uy�Aa�
](�lU������ۨD����r=V녿�P�w�1)�l[�L�6#Y�7�/I)�ƥ��O�)�&�j��TLKc��y92s�]�?5u��#���B�}�\��+�<�ɔ��k��ќ}W���uR.[0wr�4l�Xҫ����
C3v��3�Վ|�-�����x��w��pq���O,)/� !]�5��<T��];�)[7*
�m�T�!���Y��j\��̇�;�u�$͗�i�q��")����^��)�Ƿfup���:$�
���i���$Wg:AY�Y�@�ߧ��
�89B��
���p��������9>$�s� %�U��� �p���9f�7��#Lf�c&i%�E3�p)���i!�˝!S0hY%x<h}�����i:䍰�)�민�(NZv0͝�<Y�eM�= �.֜6�韴,Y�`A�팽�/j��v+�3?0����j^F�^}U�33U��e{F�ߥ�Z���ژ��xVi����@��&|�ai�/ջc}$���%�rƧ@�O���g���y��G_�Ҏj9i�y��+:�T�(Zj���r�L��� ;��Ϡ>-��(�ͬz���$����_���N��ȅH�>�>��E��wC�p��iK^��I�.�	�a�}F
o���W��F�-�'ջ
s�y2��%?�	2�sD�s�x�Y��?��a�­.sѧ&#�Q��}������󪮥 ʂ���A�X��}A�P*�@����ހKt5���%h�ֽ,��=	��2�[C�6u%�yDi�rn5�w;盖����|o�l��p'�IdJ��5	�A����hX�c:����|����������1�>��d�3f�ޭ���]�8sYfL����["A2����ẋ��%���ĵP�zXk���R�d	�Ĉ�'x��5V˻�[���j�Y�8��#�Y_%��zsij��=gg%�a��qX�E]BG/@��-ރ���,��	��_��U*�O������&A�Aw�&/il�&�ܾwS��l�a�R����2�y�$C����@"�����M��?��C����z�V� ��W>1��&Ͷ������a3����`���roQL�Th[1� ̼J���jl��f\Ȏ�XV;z�sAރfI�8a�+��N����-Q�=Z���9n�|����-r�{�A� 1�<~�Rk\�o�RM�.W��OuUG�jk���a9T��h�%�w���ێ,�2<�̉߅�hꢖw���-$^�%�JYG��[��ؠ���a,�R^�x�ﱡX��=̆Mټ�U�'��yo :r�V}oП���;�!�F�:\Z�����t�t��scp�#���H�ՉC�9�h�*�=�Rn�]Kf��]51B��K�}dl/Nn��ɞdaj�0`D�G�\���,C��
���ɐ�&i�·�ʌQ2���
ry5��c���D�,��Ȝ������N�h|�0������'_�iv1�M��oZ�<�Z����	4[s��������}+p�]���n�mN����t��(���E�pM$k��.�M��R}�w�3С����:�&
�|�+-�~X�`Z g��47��F-?�+Đ��R�aL�~�1�W�K4��@��5�O@��a㭛y5��8�/�j�S�'@��)N-MkH0&[�w��"��g���[�q�9s��<p�Q�O��@����k�~?�P�\�6��C�CGf��kd\ՙ�*��0hm����Nmw�������2��7+d����kj�����[vb����w>�&l����U��[�X''������ڭQ�j�{zy�J���h�J��Ր��@�߳��E�s��k�شo�E�@����y$5�{4De�����t^P��r���V�J2]�L���#���S��_m�g��n�2��RD�Kݐ�A������1��[\mw�竞����D��]/G(�/�4.8��_���A��Ϩ��tJ���R�l�B��0��5��Ƥ$�k��O`]  �J���w��w+n�~^���h+ۭ�',�3iS�����3[_����.G�J~-�ZH�z���U�3§k�t��� �2�/����|FӤ�Z�l�k�����'WI�Y�{��V�ۈ��p�O��
)ܹ�0sZ
��qL�Gh��2x��Ȏ��)$��F�?�4w2w<v�v��:�Y�7�H�З�|�>��Gv�Z)$�o[�;ڞI��M35�i��Y�?���Ž�˕� =�ĩ��D��#��Ђ��#��������R"�QH���v��>x�cS~�����������1�;���:��Q�o�ٖ.��Mp���;���҄���w�{�N�VV ��ͪ8�����*,���'�`
�D�"Isq>X���������Q�~�ًa�1f�>���B�G������1ElᗰRW��G}=b�[G�<y�3N��X���Mk޼hä5�L(��?�����$�:Q9��Awta��L��qXlxVHYEB    fa00    1d20w���U�$V'qƇC�.$�<����dh�k�${/k�5�b�m撲5Z��I�Ӡ�3Ń����7�g�����F7�����\�j4��F�R$��ѰgE8
xl4�mW��������y�V1�6@Q�熁NA=P��*�C*���J�ѾpS�?tdC打Y��G��xq���KFW}�.BE���PI.�~��M�{?'w��2��Λn �">ٓ;}�ܶs��Ϛ9��H�����2`ܞ����Mz�fslNj�=���=X��qL�j�_a���FW�*"t���WXb���U��]1$�r���$�Rd*�R�1d��ţ�'���d��Y��{c"[��3��5�F#R
�c9E��)�{cA��C"4�	Q#�iH�G��Y;ʄc� ��Ҧȭ�e�2/�-�6g�Z������PF]�_����p�H++��Z�9�P� ͆x�ܥ�g	�׭J=T�V ԭ�J�a]h��'��Rԓ[
��iT0գlpI��Z]Q��B����7���l���S����"	y��q�e���!��۟��s��l��Я07��o��3an���ŏ�a�&�
�:ծ�k�,V�脟�qmS�[=5���Gd�*m �#�1^76>9���Ǝ@��6�]j^1%>�D�g(E�YH. �(�j01ϸd��	<Ό>��nOٻu/]p�G�Ƹ9�s�g�RY�V���-ѫ9O�L0)�yK� (��O��I��#�B±�ֿ鄋(��7ɪ߁�A��`B��Z�W�u����$b?N���h|bƶ�_�������*Sw"�O��o==�AE�����G��W?Ly�h�����F�����q�a��Pb�A�+s���E'0�'�/BQ^�(>�����M�1�g�f٩3�*"Д����|R[�V���UK P��V&�#��G�c �~CbXc:�#ҷ�؋9��ֻPi�q'��޾RA��%!�i��U���$�_Y��n�&(sIQG��i�JL�ݩ:�8�T�I�".�K��'ސ������E���HV�=>&{8<MZ�! ˝K>mұ�3w��g�+��@@��a2�@7dOѺ�4*���ހ*�1��P�������ߎ
_�s�c�>*�	�n5� s��`�Ôǫo��6��v3�ϳ$�fuU�ns��Aw4���Dfb��������`��bJ��'�Ӈcx_Y
�����X�� �jm�֏��nO�;�hN��M`W�J�;+,�G�z(JVx����J9�(8)�z�Ҋ�MMt[�e8�d��`\���Mx�ګ��{�0f��R*d���@��
�
ʉ6'��p��Ӛ�~��Og�
~�2E�[U��%RHp�65e�T�-N0c�G��� ��+��&�1��8��7� ���2v^m:�S����Hȋ<�5�`%�Pp��.=��+��	J���}��^F8Q@({���^,�s'����&� ��u��d+�I�_6�P�뜢l�դ�龺�Z,=�;C% �����Bn�����H��q���z��7M/��h���~ڨάu�� |5�"�K뷈��	u�a�����)rC�`�������DR&u'��Q�]�m�rm׎�~�t>Z�`�&��&����D�yWە��-#����8��RcB�8\��KI����������<�6I�4cNs�O]6BKIw�'�t|gI�����ߡ��\�����Is7�
;����<�t��N�;�`����r(���m8��Vg�~5�ǳ.�"��޹���LAø�u���6=�͛Z΋&"�5@c�H�~2{�]�3<Sݼo��7v���ኺ�q��) �jdk�%ו�I��a[Ű�_�$#5u���̷����h��4noV�j���%���
��ω�h�!�r5Pk�,?Ih����9;��,a��l`��w/��*�(�#8���i�.����oM��
�!��J��ńqD�/L,ZD�6֮��7��W��Ɛo��l�7�t�� �	��mx$�9�iM$ �*��H�#����0ޟ`-G_���u�..�ĉmډb��U�LK"`"!·<3^֊�+�Ȟ{�5ڹ�C�?�[�~+����u;ob�ˁ(!ҷ.a_�@��g�J�L��]��Q�I to��a��B;M�W��(���T���B�/�_t(�]��w��`�(��k�xCfX+��<�h��r�=�n���D8p�OXy��W����4��;� ���_D<5�DS���]����\�fء���fA�L�6��i9������:P���mR~�nm.m |�e�G�f]�Z�?��N����6/�#|��|�f�	��h$r�(}�ew�P�,��*�]P�P`��迨�[�k���C�W� ��H����c?S���Ս�]�##Y�$S^ �ɛ���]�&5�bפ*2RQ����̠*�16g�L�S����N���%n�����S��+��Ϸ�\�����<^@^�X�D���2�c�a��;����	�&_�"j�U���pZ�Ll�{u��K�P	� �p�j\���fY� ��-..ƾ�]�ڳ�D�����ϛ��餶��������xb�KCc�*s0�ƃ��\�cM7[ݴv�t��
���DkwNVf�t�{�V=8Ϲ������l��:�'dDh �� �'�Z�É#<�2����<�;�BՎ�Ӄ��Q��P������0z�+ �1i�A5���5�rF��H�U���k��X���!��!���T�C�H�Ɣ?�A㐳��ۙA9�M��.��ѳ>�W�,3���(��XLq~�&:�0���?1���������:��r��V.15:����嶂*�UhHM�����L�����bk%W3G�Q�������e�B<|j��N���4�^d����m�jj�֫@[����<��N�x~XG튕3�	�x��>�:���B�*�	���u�,c�V�\��h��U��n��^�����@�]�-T\0?e��S������^�vs��a�r��x�5�	S\�5��q�0�^,�GGf�'
K7rE����o�
�#�$_ �nv��ʺ��p
��It8h�,bs]�f��;�C2p�jaV�	L�����������(�wѳA���+�e�����-k��)9�_O��{�:��}?a��x�ю<��|1e廇�)D"��x��/����la��v�A��L���U�9z+qdl���XyߋSBë��:N��(X�q�A�"^��$��aX���,w��N�������_�-�e䛍!_�)������\-��;U�l��z�<$QJY13"컹��sX{���	t��2�iV�:�Q�-��Lߨax\=r�$!�� fPs�?�4b���\ỷ`(�uא�k����@GHcl�6����s�v�fTq��*mTڵ��v�-D��Q��g4���P�O��,�����'���!ɡA���k�41
j5^�"��Z�M"c?h�6�(��4[ف��b�XK5}kR93s�����\*{QM�D�=����+mnb����NV���6��'��!����e������/�Ϟ��U6C��DmouA��E�*�M�?J���e�?���z6�aY�6����˴C*������~�I���gX�qt��`��R�I�g&��;��;�	�r ��>y�l9L�>_�:М�F�Q��8S�NÀ��tl}xJ�gu-X�LYW}���rtٲdL�4��8ľ}��t�3�����u�F���ۗI��{�	J�aKW*�M4���H6��!�J�̡!�1�'z=� K�XBk��*���d��s�����DS�7��5�:p9wyp�A�𦫁Mv�D����VZ��.<�~���Q��G|꯰��K?�M�����$ix��_�9��Cpؕ�]9���F���`��J����ZT�9Po�����ݷh�c�I����puycÃ�)�]�}���)�Z!%E�-@�)9��\T��f���	�]���;=NW� -�"�Ke#1{�\��'��X!p߼^�pP4'�R����(��A�,�>N��5��?"�`N�*���]T?�ǹ���H��F�I��x
�x&n�Wf���w&��@4�A{��&�;�p��B;���sۮq
��l\�b9
�PKr�Г�y}�e�:��2:Ռo��� �9-�]���ϰ��+=������?N���h�����o ǃt�����e�D���b��ۘ�O���H�,dR�����F��o�b<<���(�z�HT܅�M�Y�D�W'�)k�Hm�Db�fq+c�9�?�3v_�s1��7͹�C�M�|;z�:�	l�!ݲ�,�T1+��i�tn�E�Tx��Ry�$(c-�fw�פH5���)}�Lx�R
��U�Dqr���E��;��e�G�c�F��"q�F�I�b�_ ��t�yЏ����)d������XYC��"�g���ﰪ84�ٴP���yd�������;�U�[�h�IB_���$� �pQ��h��>;A��wkln}��/>��jv\�b���s^6
��>AW9Jt0�#��g�����;Lw�u� +�����uh�,s��h��6:�L����|�R�=�I�v�;�l��,�@�"�k�cq뉝���g��� �?�uJ��A�1i-�wU��Y)���q��?$�5�<VOL����U�SQ���/7-���}"���E�<�a��yB�������̚��;���/�z7TQD�m3rTXUĲ���nG�����#K7�,W.k�`���E�pv��A>0
H����/9��p �Ґ��đ*�x\N�L��w��?����s�$8�1����%9��'0�Y�Q@�O�x�1�V�?�+���}Q��Q#���JtB~�$�F@+����W���e�p/�3.?�ʂT0DR���!��Bݛe.���V�����M|w�(h�V�)C��d�����6���}��<�O���G8sn�ztN&,o��g�`�Z8��ѩ�紡���N��%
����oP�}/�s!��?,wf���%����Q����蠴���Puepe���dw�� W'e¶(�s�#�����p�3��㇙wdM���?o}��gu���5C\:\���;k�kg��;D��L,�7=N��ES�~?aB֤8� 3�+�Y��o3x{/�	C����;�1_+{-�Sr����c�B�V鑾.LiGC)|�=��m`������ݦ���Z�|?����������p�{�Gܢ8t�u[L"��a>�<��b���"�W�����
��8ff��؂��Tq�zR�t~��0Y���	uJH�u%s7�[���?:a�*�d�'-s�<�cA���]i��Q'QVŹH��rQ����J�ʽ�۵FMI�Q����g/4�iM9��J����J���At���i$!}�����u�V/����yEQ=ӝN��m���=���g��y����I�؇�.�|D���d��Ëg��?���=�,����:ۋ��G\��$��bQ]��h#�I�x��{hkS���5q��Vɩd��)r��n-]1��5�9N���p��-z�����=x���]#א�2kl!F-=
���L��^�G%����]9����'�����=ٷSd��q2p�+�*����IA�c_�xJ�a+�<�D�ۓ�`�uc^�h�A��������Ov����8�ֶ��u�5]���l �QK�m��}>�<x��ՙ8���J���p��hvV�S��-�3��Lhga�`��Z�͢�t�π$a`��M6<����oQ���4v��<Y���x(_�+zkS�j��D;���Yh���z�0a^��c��{˚el��aa6�'I�K�WM�	ȧ�k�U���u�8Im��ܵ�!�,�5�ܹ2(8S*�p���%�Wg���DWMC�&��9T�Ca��d|��G7��*UH�4R5o����fHmh�L�2���ԅX���E�{K`b!o�Yy[HƼ����0����㪌R��^�niF�j���껓,)�*� |?���+�Z8�]P���ε�YBrޒ�<$�D���K���7��.p�[f?o��L[�8�+�y��U��=��0�Mo�Sa�i\���+g,(�z��B��&FǠ��D��Hk��2x�L�<���V����1�'�~��B���0n���P�;���@�Z���/jϻF�>��\�lr�:��Z�"������*�aP|�H��'X���hS�KF.�����A��g�qu���]��טN���D.KǴ��ӄ9����J��B���Sfmom�~ r���n�������C��d�͘�0��	����+S$`婵:`�<�;X�a�;��
*��
,6�3{f�K��Q���0mr�&Ԓڈ�.r��B��]Yǟq��nqMw�S8��L5��^�'Z[��J�u�3�zo���-V%~���Mɧ����E9j��|�ثu������ȍ�@e���dY��W�g�u>S���\��f'�?R&�"�&y���_�z��8��%���>c6Y�4ݨ�Z�Bi��%
�U����Ǥ���S�KJg�%\TI�w�����f�%�vEe�������]�K�d���ӓ��k�Z�����}aE?=n��R�0Y�۹�����"iH��L���ңp����^��9��Q�������ܾ�����=eI��ⲕ>rn*.��w�[���z>��ZQ����0�FK�m�)x�v,�q��O�J�61vi�c����4~v^�����R�b�J�Z��&*�/�7�aBν
{����h����&J$�{D4��i�&�bל$�}�'d��� D��޳�XC�1�)y��͸�wD"�|��F`A���ZC8K�;�:x���l'�<z5F�a�t���Jt��%�V��!e����WIl�6\�R����}je�=��k��4~p�v)�YO2�ϋ�~3� 	��07�5�0���C�sի^HU�d�%-"�ew�oL9�Z�ٞ�ޏ�K!�ߗKςĈ("Epbi�uW��a������TlF��
w�:YRj��JY�E�%�N+0�]�	����#u����UG�c��k<��e�qk�I~S�����:5������=`��������c�Q�|�����O#5�������쐙�nG[�dR����t�R��q�>"
���K:�p���щ�x�}@x7��*��G���;������'��Nj��0;sړl9P��Q��:0��)��.�]&Ѥo/k��!A,"%�~���O%�2*���>�T�N��}�.XlxVHYEB    fa00    1e20*H��.�����2�.��::��W�W1�֡
{��Cnf�=$�o��q�/�2�a�i�-���{b#�k��n�S(�����j���z>��f�ɻ$�@�GŔ�e�#�3O5ȓ=�8����!�� ��GP���G=�&�F�i��0b�; ���nBΜ��L��_JÎvP\w�j��|ј�ݛ�Қ[�lw��3�{!(�}�up����F 	ؔ�D� �&���{���6o���{����\C/���j�;�2sa���iȲ��!�ȿ)�b���b�?J;2C`�3xGI�������Q����Eb'�su �ه�J��{���'׼�̴*�E���2��tJ�
c=P7~>��oHe�K�9z�[@����X��A���0v���P�9���6���$�~^���GO�M^���	�##2/g�$6xP��m�{c%"�T�؎/^6v��يr�w�)��-jC(�`|vxp�S�ؖC�F���������n�U=�N��D��c)Ay?��?�����X^�ޔ|��?ϐ������y�a���V�Ř������_��a�����&9D	���σ%��'p~+{J `xGVI��c�����Z�t�n7�n��%�M�-L������v��ȸ�ZD�%��+��]�>=�P���1�άF�c���I� ut/�C�4$� �
��R�F���o�B�����ԟg�%��Q����xͬ��],��Y�H��ۿ�R�{)�1��>,���q��bԃ���nb6\�^+Q
�x pN��=ȺD]�����s6��>OM�aʡ},�_��E���Z�穎�mL��(��}#J���3�KplYԣ��%PS�d��!z{&�?K�i��U6i0�f�"5L?�8�d�>�U����5�D��t���I��wE��~)5s�hί7ʼ�.��r��Uգ�#�m+�>׭��J�ػ�T��(TW�v��Hw�VY��V0[�RCju�M=v�; y�3e�T�K,r�,eg����:�zq�#��%X�7��	i�2�ɟ;ӯy ��O@�i�u|��-�ܠ#�W�}X����.J&H� �*~����G�4��WD���]��i\�U���,ͩL��{�o�tP(��7�ﬠj_����A]*��w!�
�G�i)�^)y�2���,.��G.X�Et�x4�a,,cDQ���^�o�nH�%��s{�Tϒڛ�*��$GF�B��K��xNu#1C�z'Ҭ
���$��Q�|o�H�06�N�t؆)"�Ͷ��R��B���!)�N�v������WX$~��wj1�ٟDR����eh�R͙T�Na��,.R��^?1��y����%9D#=��;��q_�x�J-ɉP���r3q2]�Y,Ұ�`6Cr՜t���go ���C�A������MH��M���<�f�reC\��II:�J����3𧦦����w����T/E�i
x ��ᄨ{�&^��ls|vP�o�q�R?�����:�	G6߉�gI>tu�}z�u-����D=E��?�yys�у<�<(!�g��I�L�fz�Y��gw)��R��U��*��W�'�G ��uҽx�$�6��N[����)Ѷ��7yi���uas�ɱcZ�$�~oԥ���"(�o��8Z�?�G5�L�Q�L5�m � '��O�HN���u�a~�D�P���`*ǹ���hr@�X��E�ѐ&�<6�A��WV�vݵ��e>''d��%�A��}#S>�\;w�9j���ԓ�_�>�*�k�1���׃�1�s��:g0(�i(F�*��ח7���m����q�ܭ�p�%��.V��S��:��b)� d�z]�jD�l0�+�]����h�9u��11�Gqǻ��hѤ�8Z��!N�"��f-�w6T2-��#H���E-s��)x>�[?����FΙR��HX���=���k�L���iw�SÁ�C���Fh�kБ��el)��G
�{y����*p��֨*�f)�������;W'j��6E�>�!�F �p;dū�Љ5i��L|��N�M�0�Ƣ�/}��Eܸ�������˭�D�ꑬ�o�#iP|�� �i���I�Ck߸����J _�4���0ڄ�O���Ke�ZB�e�3�2���*u�O�cJ�^��"`S:b�>@��:�!�]�C�hcwļAϠ��o���-�iN����A�t�@L=cs�6|l|�՝˰i�x�p��q�'f�F�E����^'�§��{$���z3�#t���~,�)�uSb�����j]i�͋��n������w7/��B�SU��hl�#��|�U��E����Y�)�%c��U��H )ű7ZڔY�.��.O�b�|.+\��͋��2A����@����xf��*:��B����!�0����C�dl�f�<G����c�kЧ���S
�567N$����1�����l����ƀ������5�����܀��Ͻċ�qɋ��osT�x��$c"Q1�Ftu��7�5�ta�.@��f������_-~!��r8n{����=4~g��l�Yfa)�e/9w�=@\u���������Gb��^o�Xģ�c�v_Mq�`����xus���<�A��evE�_���(/��/х�ӏ�:vm����IT�⶝r�҅0��2,[�Θ%i��T�Ryq릁KǦ�ç��K����t�5�n曄�:�I��p*�������+�2k�=��|Wįy[�
�*�mr��e�+(�4�hY�o:X��o;�m�� �=Ѵsu��S(�TSbL�a\�;��VDv�,������p��oO��(b����7�j)�$��	C����6%GM���+?n�/����N0Ӻ�8���[���{��r��;�&�ͫ��y{b���L% ��s��|�;vYGf��(^Q�*Yo��/UE�9jT'�-U�N�۔��~Y6�����{�jG���V���+� ����zx���f~7ca���ǟg��Q����d�: ���y'���0����<p���qfˋ��8c0��M��i�a������3	��>�)[���';�L���컿X)n������R����m��O(Gh��͏ᨷ�g<s�ͺ������T\�:�S�BQD�Чxx[�7p`7x�b6Z��_�_g�q�0Iщ�T�z�No U�5.'p��Z)�JQ�w��k$hl���a\q��M�)�%a���ٲ�S�n��z���I��FW��.�-��)b�-�� ���XX��皗��j��	}�۟�6�݇b�QIC�^D5�v#��<�A���KwA�	\��!=;@�D�rz�+H@x,��"}^��{�-��Ǻ��c��g�y �*���+���HGq�2��^82�y0�/[�.��"���n.ӊ�k+�b4�yKx���2V��<��=��� �r�=�ң�wT������fCS��
Y�^����?�I�s�F�~�q��ק#��B��B)���,��k���\��\���6�� ��Y�K���խCjZ�:�g>t�]���hckM� �H!�#*�{�M�	r���qSއ�:������$z�D.Q�sQ������]v��=��h���3�U��X��ŗy��Ǥ�%�š�}=�����y��wa?�Ej���o] ��,pJda�~Yw��vd䯞psr'���!�%2?��J��QA �L�a��<��h�;߫{��)����l�Br�)�~����g��e��ds%w��Z�Xy�Su�� ���c2%q���0eX�s4��&��yI~����Z&ɮ���i�_E�gò���Z�k�tZ��HL�m��+m��7]Bo��*Ja�0څ|K��«�x3F��OX=O��,+G=L�j��T90�?2�B]	�ȍn�"l?����F쥸;V�J���`��e� e}��	��xy�/V0��߶� �3."��G����e�9~�!�Wݾ���uX@ V�6��*f-�]�c��s�vr%�+��K�7�:;�:� �3�z�\lc�ok1����4H��MT��8�E�~�Z6&hj�NH�c28I��\�4痐��uh�7Ea�������!���~ 8l	�	�߈vdi�uV�:<��]�O�6⣄�yo�Ϟ��50\$��FY�6���ĉ�(C���là��5X��K��O�P�g�.�tC���H���]��R�lg�����ś������Ww@K��:YjԊ�1&e��2�Q&S�V	�ځ�K��E����b���i]��g�2VR��#Y�8���#a�_1�6x@=�$ݷ4���Kױ�����Ƚ����׿NS�Eu����d�ǽv���l�3���T�����B}B��x�D�Ǧ�Hq��v�r��M�W�j��]H�XfT��㣺=�p�����߇�xkf��20r�܅ɂ*������̔��zn-���e��2���,��@ ���i��ሬJ��s"�v I"�aER�_��јceU�RV�;cP�D� fc�9�5jiȔ�l��C�L8���U_�mM�����l�D����t��p��ݟ��H�ԁҰ?#K�-��5 cY����Hy�?y������֝~Rg5�.�<�pEKyCi����/*k�0���;��ѣPF�r�S�˦�&�D�x�r")%;��eU�E'��*r&`RG��^~�삃Ũ��Ӽ���h�>N:"����Lt�u�}�m��=BS*�D�`�*0��2���:Z�G�3a3��H {MSԈr%/.K�h�b�Y�"��SȢ��u��{��J�G����e@�i�T H�r_���e�c��Rb��܆��j+�0��4ΠѺ? ���M�� ��\��X��H5HB�)����R��}�?�N�wy���N}1v���8�����%�{�.���ש�f9h��b]���:����{���v3�6�Z2�n[[fZ妢�[�ދ/�KdV�	Q��[��0Y���qaV')p ��5�P��O��<{?��VQ4Nn�")^��D�0nŔ�o�#c^�k_��u:޹NWnR~�}IV��d1n��|�/ֿ�C�xU1�7�x΁�Sf�hH�p
��3��4}�1�)�ྱ��J_������}~L��V�~k�������'��O� ���R�I���T�ì+ۀ[�"��{���[�9N����GOC:�m�E\6w�"_����Pl�����r!k��(�B�f^�Ȝ��T�ߛ6 ڸǋ}��"\�ɩ)Q�\h��o��b���g�ZoYԢ��Bv� Z%�(�x~X���N��͗Q�]5�;$	�BB�q�+y-�G��=J߻�I�(f�v���4�%���]<��(>���Q�p#G��a�;$D�@|��k�
H8�lD$7�l8*��oǘ,��{����0\!L\V�K?)�����a�}u.�e����pٴ%��o����$��	8c(S_� �����
��$�O&CL��t_Ns�ƈ7��l��ڋM���ZS�"��u��z�}F�(�&��su��9�@g�e>��0k���M�Yl�~Yo���$ۘ�Hk}T�n�����bU�P\�qf(.�N����b�ǋm�A?Z0D��+1�	�VB����D��ĸ/{��/t�.+�y��26�i�0Ϙ����� �|SlC��lx�������P �r1{ �`��{�A�����r���B�L���$z�r���]U^-�]�3[,������4�_��r�*���j����(N�IO�k�-���Cu<����:�\J���QF�ٳ��H-�s!-������fcz0�Z~m��؃��^��j¿�¦�.�b���õ�l�ӡ�m9IC�%���)��]iT�A�e����P�=�&��^�U�Đ���yq̎=Q�T)�29p�u��\��T�k1&�u�X1P���<曧��vv@��� :�0�Z��I�lF����4En�Uu�z�����7����N�ynf��e�s���(f�o5dJx�Ű���f���}�\����6�t�=e��`��e�z�b�j�Z�MK�'�O��	�%� @�o��c �/�u�E����b^������I!BJ1����A4�n_4�ᖳ�;�+2�1왓��-�?�"��$ׇ�r�Y�#�3{�Y��(e��n0��&5j��Ɩ�5=�}�����q�9/���E�Q�:N~Ͷ<�(����P$T�h��*�
ܺ*��]����c���y{:y�z�N���}n
�W3��ϑYq_�@c��3����*@�����Ɔ	tw��A������,�#`@��p|)x�%^H.����-"��в�l|�N�1v�j9_�]Ą����~��.���[��-�2��ր�����&�S��xG>���|3� qnܫ�y�/� #J���F�,\%= ��|*��K�O���:ע���Yޔ/@1���IB4�%�% WN����>�&MyӴ��H�j�= ��@�sL
�w:v<�L����>�X�u�H0�h$µ[<���4-WHނ�~=B$j���$���Z���k���x2�̙�r�*nꚆu���C��R���ט/�Z�1�NF�|@�H�%:�ϸ�1����`�%��z��A�]/Z�yS�*.4&��L��_�J�݅�SVL��>l���	1��|zwvÜ��}�j�.��?��+zM/ Y�x"�u�����%�1'K��*ݧ�9��czf�3�GiQ�'Vor{4<�!�y���I�=6�F�lc��~=P���(P�AF�!�k۳l�Ж����+f����.1n;�4��X�B�*EE������U̒��s�U=p�q9�p�������Փ�c�o��1?�1�5��G��S]�A�Ľ#�}��[&]Q3kO{)��|�S?��(U�<��ey�^N!� �h���n�B	�|����)��aK7�z?aK��Y����G�h�Nz�C���Vȝ%լ����)��WQ��;=#�<��
����<�)��5�fnQr���ܸ��
p�Z\�Z�^�loBk*\\ƓI�V�ޑOcIP�3�?�7�)�Y���Z��}ST݌�B�%fE��S^��̕��ٖe���KXU蹅q�d�r��Ȩ�Q��}ڷ�����aDk��R���(:0�27a�]?��B��"��� ����go}�T#��+��|�m���de����ԥ���>�Y�V���=��b���"\�S#&[�x���\��n�5�J:�=�Ba|T���(�ݏ/V����Zl��W����E��&��&�<!��>b^�fo���x[o:;�H�����Y�(���ρ��Ğ²���⾌R�Fl~n�q�FU������8ܺ���9��X�ݯ�1FѶ1?UrZ���v��$Z衬��_yL�����&�z�;宯Ad�6���ס��/�HA��=d�D��Ku�J�¦� �Gf�`�W70���li�'զ�M�d���g^Q.��w� ���kHƕ�2�A/�UQa�_���ps�=���᣹^bP��'��3�&�#���V#����N��h�oQ:�-�a�9J6#��j\�,_.�XlxVHYEB    fa00    1e50�(��-ĝI���a�/m#�L][�Y��kqx
�������{�C�8s~�0θA{�f��q;4���Űŕ)̾�~����׼�U,��Rj��Zz��]�t �t?�Ss��vS��!Z&�kd�$]�J��l�ѐ�*���W�IZ'�=>�m�־���W+�쐰G��9c�:ؠ�M�|�,�hw�~��~8,�.����-�&��9�3�8
/5ЉZ �`��/¼ܮ��^�Q{i[�LP�Z�
�.��=�W�E0(z���re��;^iR��s�֖N)9���:k��J��a���q�I���%�����C�A�V�-��T����=?��� �$�xg���O��v�F��1C�@h���õR��������9�.��ri��%���Ѭ1�K��w�vn�p�ř����"��:�րb�^�����3��P�~�A��1�v릪~%�W�Z��)�A	��gb�Gɞ�R�4��WI��}d�I- ���pwV�sv�/{_�Nk�¢���T1%�Dd�A�Eq>���J���n�ڙ�/?07*^8e��x���G�<
(-]�����R3���5����@�$�-1�:�1\�D#��jk<���M�|��۝��ӺÂ�=�Ֆ����?���H�B[��ށ=,��:w>CR8 y͊�o2�(�W�Pa2X%[��&��&��@c��quVf��(�܊���c�x��iqo�c��A|zL���,Ĥ��H��I�P~�+���7��V~?�l���c0+<��᝜��EZ�~
��E�� ţ5��HB)&���t>75�I�Α�ញCؒA�7�Y�Ʉ9��:Y�L*�����`�B�t�PMΏ�!���Ǘp{�DXf��ggE�����ٛp%�-<�k1�(��ZOҾ�Z6Q	Wnw8�7PF���% �R�Ϥl'�L��9f��5�T/_�F>�`��5����[wf�:�Z�P	n/
<�t]��8����,�aA��k�yc�)���n��O?��sGYq*�:�tc�$?��J��;�v>*I��ɥ�o"���hAx�1H c�"^�H�-Z�UD���V���BNւr� �]rD���$)Ia�/͔��|^^��k���2`Rh.|~�zc�爥%hm��ឡ�)�Ws��ܻ�Kb&�>4���;�.��|}lN��M 5*?h��xI��c��]O����Jj��r6���IJ�'��?�����MA0wYGe"�ՖL�7�צG��^;j�T�F�s�6���ȊP��	+���I��P��R��²Y�&B�n���&�^4�7H2jt8�RYE}z�3[H'������w�`e��h9ci��;k����*��\'���?ލ�석^�����Q]���+p9-*`�tp�	zE�7�vR�nibןwo0m;%��M7ݼ|�'��=?ǭ�Y�E�G}�QT�3	��:��)̱2@�st�ܜ�wV`]Ù%�窔�D>��vd�z�k��{'%l4�,-9\~R��jFL�v���a�M���	5(1 o.۬�o���s^�y7�����dӍco�;CV���ˋx[�{�a���]�|�Y�N��nE����  ��lB���	��ʡ��Ƴa���2��1G��8C<);I��@l�RL�F(��h�|��Jj��@���2���z�� ���!L�}8������nn�Qb�;g�)y� ���Q�{k�r�%�E��Z��$H�
�.F����C�|����L�Պ��$
ſ+u����0jA�n��[8�g��	��s#U����c�����ṓ��r�]��N��v��c L(���	�=+2�(b�y���O�"��K�K�X��_"D���K��ZZ�ST$A�ގ�O��hY-@nb����!��������u��սq7o��F�7�'sf������>�8?3���=��������-�`�"�jc�4�n�Lc�l߆�O�%_�a+���fKPV��b���	w���ª�w�/�G��d`�}>֮�9������?�2E�f��3�İ;6��FDAș����jV^�������*ףMs�q0nyw��P���$��ηw���EY�N���2��P�^���;[�ǿY�=������٪6�橃h5�1�"����$8�Q�#�Y�_�2��/F�X)Ark�a�:!oХ_�4��̐�J�y.��F����ƍ�z�Z 6,����=�J���熍RE֟�7�2����+�.w�+
��[�^T*�n	�g#��N?��f�0�R�����:g��3�igR�����af٠���ф��_��aV��|\����s�P�js�h��
�c�d�P�д �j��7��8�B����U!O��}o.�vD�Q�N��/�s����=���I�Dp�d�|��'�����I�?Cw�L�<�S8̇t���^>��#�01��sz�jRxp0c/읳R?b�N��lm��ćmf�f'I4����\-ƪx%�tF�n�2N"��IB��J�P\���� �u�5@�i)��q�ͭ;_j��OG��rv�i����i�GSI�(��E�n���f����d���S[d�I�rRXKN[��]'�0�	��ä�D�f�{�n�a��QKL}�Q9�1����;y%{�p���uE����8�!���,�C��87^y�vј,�_@��մ�7L� 3�ͨ?��wG�����$$�c���PX��?��$y��!E�[�i��$0�y�a��f��� ������^�+(�9� <�Eʸ}�\��7����+�c����x~<>�Q�g�(�g\s;b9%�4v����$}�� F|A�,XmF�+2��i�̎�Y��k�@�[�h(��~iv:~vh-�V�����r�q�� ɼXD��;�ri�y����nU��x��w��S\���.�q�}��+�������I؇n��%,S%^O*+@��:�wZ�>kq1'Kq�%�*y2�k��,T��ݍ_�j��NYs�����&��){L��[J�n����߳��~ڲh��ۋ��V�Y,17���՗��UC/��t��D+{�%�s�<8�U��$��4�`i�w���f/�nu\ۂȏ&aH~�M$�N4���@��C�=DJVci��a�l���ol�(o��g���s�-��F�t~[�v?�#v�b}�l��&u�ˣk��BM��y8b��Q�k�*��_���n�O��������Y��fF^]mg���|I 4����b���s|ʕ�w�@�β\D1oT9���+��8��d�X��*{	e��b���:�D�Z�m�� *u���� ��<���94�x}�r�Z�:��<}���[;@�d712W�\�V���|�ɭ�!�u���:�,�NB�y�����R�,��m_�~^fJ�.�%y�N�daF��@(��U�J.=nS���I��6��\e4�J��ZNð��XNfEy�E·K5o��:L�#�<V[�b��.�( e�JV�u?^Zf����}�D�?wqIz�C�鎡�-�CB6�����^}�0���_JY�1}D�U|/��f����a㈩��o��]��$4��=a�<�F���<�yX��YQ�:#��'&��`�z
�9��߮��hG�Z�&D�1�:�h�}���7d|�Ȥ�q��֬ 	�bS3a$��d��Խ���{�U��?����ĳ���;r����d#�Q�O-�wQ��cO	��X�1�$�� ӳ��N��(u���o$��(�卭�8�}P��S$�0\0u�*5�]��S�!�R�}�M�f�6~l`�Ka2��W�Z�ęL���ڷ�]���g�rG�R�u���<��|��1Ryh_T�?�kZ�r���W�g���t��U���@��L,[����JbZ�zK��S�F���=�@��y�6�1<��%�#�:s�HW�;ڻ�0s;|���m�׆��	U������,�ϒ��}3��.Y�<d�M8{���C�g���Z��4K�2�ݓo&�S�?�ї3.��,O���Wc�!��ɧO���'���>o�+u�%�5L s�]��3)^W��\1�"c��n��s@�UP�n�U�9}	?#w�;����� [���8��6R��v���3/B�0��EU������.~�>jB����d5&���~� ��Y�4h?	���a~��GR�:�&�+a8��u���̀�XK�U����
9>��V��!�cN��
��}���b6�.H����t䰟�7}{���QL[j9�(�����Y��#-UC�_�S�(S $�G<�An���`F;u��xAC=�t:UĝRH�ո�ӒRo�߄�;J��Z�3h ��9w�z"��`�+?��.�j��}�.:
FBC�?�9a�XҮ%��!eQ��
h�{,'�/��5���*�jׅ�	���c��?e�~�C�4(5��̂�~ӯF��6	��5q8H��Q�I��vŘ���w�2�پh��)>+}W��h�_��
���`��a7�c��h&�~.��A�e.R�"�M���^5'ƒjͿEź��ԁ`>N@0�=��n\3(D�'�:d��VoJ�Z-W@�Ҏ�S�*c�{nU�A�o��+�
z��D�{T�`� m��ɷ���:�J���p�/�Yr��K\OY���t%s�en'N�@E�kD���됩�xJw����ےC��Y�W��ud,���:��=�:lH�e��0ǽqC1:�-}�~~�P���-��Q��ĘR{P�Eoϋ���H,�e�0�7Q�u%��hG#w��qtA����\ P��BbZ5�V�D?y��5��|���9܏��) o����=��ݖ4�,�!4�p�3�4�؋<]Ѷ�����C{l��"Χ�I}����dE�� m��� k3m�΁�)���(���g�8����}�p�~�=v���m�U��UD?��[ ���9�`<!mwW������k�Y��4x1 B�~�=�	�>y�>�#���G�e�\��:��]���@+���0z(�;�c�/~��հ	�Ц�w�N���YId��(U�>j!k�Z@e�<�K\���Cf<��*���CO�̩I�;��u�ԝ���3�i�Z�"Ɗ��V�nՖ�Q��Dl9j �w�$�5E�+k�åB������'V�&V�x����g��C�)$[��;�Z��+��MQBUȖվX݆����c��y!c��-�|i֩� N�VC5\��ϟ���� 9�Q����v�#�F�#a��7*�R���Y�9(�T��������$�M�(�.��hG9}ie`�q� ��n?8! �/��������4�l���N�#�G���G-"Yי�*^���761�jYL��6���{������81s	�\�iQja��(:e!�ߖA��a�(���|\�z�u��u-�o�������᧒��2���<,W\]�k�1)J"Cf�|k|�|L���|�c"�1����iO����<1;��C�8��I0��*��Ê�hChW�Y.)�鐿��w��7N�@_�5�H��U?�h�pU�]e�"4wθ@P�M�*��.�`c���(T_W�W���l��?T�LBu�"V�T���'Ehx����\�:����;�1ɅꙄ3U��d���eO���rV>���.�kJ���:�aY���,�̰�Zy;���!�|VQUM�{���L�z��𢻟)5.i5r�OM|��d�g�+���6&�D}C�g�P��M�ᢷF��=7��5?��ʰK ��F(��;s�<�t�[4��ø� T�B�t�o��tx�vi��Ͼ&��d<��H��C7���~��_'J{*6�5�}�PFv��6�-v`��>%��@�R���B��Je�fQl�$��������q��*V�*�O���ELݭQ�X�c(`��k#����!�;g�?����19q��42	X&�7j>�s<濌Bbv��WXW�Jv�z����O��A��zs*Q#�'�\���e������*OY�=�`bR��	�i���X�����bMJ�i�:�-��q�t)EJ��<|(�W%q@�]Dd�����2��f@��N�Ӄ��r3�k����/ҋ9��p�ؔ�;zk��dؐᵇ�<D{�ByxGg��)�l� �1;�����<�y?�@H��S�4+���ٍK6�ӑ>�H�_����x�7Dj�zt�wI,���w U�ב�j���J���L���3�K{s,�#��ܳ Z�g�1_%,���2��dG�yZh`�w��0�Kޔ�M��PG���X%�Π�����#&j��1�
���"��u���!��=R��]��g�/^K�����������]��R���:�SY8�<�z���~3.ţ�H�D���{�OM!�G��N������{�r[�T&��y'��+i�z�����;;���g�1@(:��V����ܝ�S�[��HI�g�X��N}�1Xq��6�����r��k�DV �s�;j����[q�֐-�ud��A�li�g�4��J�	�%�4���I�fň���v��E7���T���5���j�!fW�O��7��0��?9�FW���-�p�:~��֗f��e�
3��0�]�)�0������~���	�q��Z=!6��s���1�6Gp�����RJ�� Rk}Js����a�|I��M�fX�%ȣ��w�3�_�+��7_^_��
E��O��P�|M�t,� h��'n��dv��^��DW���&���3��Be�f����h1�{b?Y�����R%��X����yX\9��L�s�~�-\mx�1��Y �.4Obԗ���%��#�VJ>ao6�S)|	�xL5(�T��{sŗ턁��ǽ.�/�@�s2W�v�^V���w�o��Rȑ�}������t��(���䓤ϰU�z6�͝�K����H��`'W&Kh%�-q9�����h����YǮV���EJn�П�/d�]\�H�S����&�CTYfō��W�Q�)R�WYW��f�\��Dk���$c> N�^�P���w ��L�ʧ�}��yL![�|�si�,��h�q
f6f�G��Բy3T5~؂^���ʀ,��H����L ����fϸ��E��$��wBz�Gf�b�A��7� d���5��B�ݔ�R�$<�=YЗ�V���Y�=$p	� �S|7U�H���^a!��jq�p�h�P���8[���Vr�1�B
�{|���@1��AXN����:�/]%��|��?�g�ʄ*^�\�Ҹ�3D���PSo:���s�i����V�'&�[@�� �A��n��'�S�`�o��n��{��;�+U�Y�8�K#���D �%�42KF�h�}�Z�Х*�!նaJEB�MJ�����:zE��dN$`�A�D1��or�(�U;}R�@�^�Kub���wtsA��1*�(~D|
XH<(��kҸ�F��׳qB5tw�_cQƸ��D�AS�D���{zeώ�͋0NZ��\؞B���LG-�B������7lec@�:�FRs$��A�
�E�Pc�P/�-^#�����e�����I�~�b���|p
�C���❬�F�́��{�>��pq3��"$c`�Z=p�F�!��LI5��+lo���b?��}�����v�$XlxVHYEB    fa00    1da0{�y��l�3����s�W;��[���[_f"]dnǾ�A���>ȍ?�sy�zs���R��HOM�����~�&��_%ܵu7ٽ�|����3��͉��'���N���׷Z�mO��@��m ��I	�^H� �*1���������4)2��_��^jc8E��۞�ys�+�𕻟�	��� r'Bd�v�3~a۪�.��)�;��!���m�2=pkU!��yvJ��E�� �������v���T%��M���!q�A��5��=Ԣ��*��_�X���ٲ�8S��e�Ri&h��OK#,&�-�K�m��?��y�� ��=�H�+�!�����	�@�%��f]�:���]�d����Q��f>�n�V��%S�����#�<8�2wnp�]'s��]��/�lh7��_�}>RV$U�䆵$�`�-�v��y<�`��L=s7�q��כ��4þ�T���{�:�o';E�!���`Cץ޻WQrܝ݊MWM� ���c���A���/XG �b�^vԭ�
�`[�Ą�<&F�����N�X�`[ʶh��tv�R�)F�xv*�	�c�,ptȲ��͌ۗ� ���o�׳�I{y���iu�e˸#u޻� ����<x��mӚ�R�^+����� �������WJ`��v��[��-ը��]�$���c�`�.�bz���z���Ϗ��sq���ܚ�2�~�?�j�&DN$�X����n�y�K�@��5���֧��Ct�"0��S�l�R�c������4�'IFai��8�4���o�ƀ��N����Y��Rʺ�qWⶍ��U�Ȉ�\�xw�{���Y&,}��]
����V���i���Jd=$#��e�TGu�� U�u;�$"zܺ�v<s��M�>iM�a�47�t��,7������}�$,���w���I@�`Lܜ ���M��sڲ�v1�}Az�!y�cUz�&�V51}�����Ѝ�P~6�L`m^MF�0��9��m�#�Z��F\q�������M�SUtt�ҧ]���S��g��Uo@�����f
�C�![�� �gI�a88оce2��ڹ�m���P("���c�!�� '���.O�?�ޑ���jrO=�4w�^j��X"��x./�iOqO8�9�"kkUwV���Y'|����,i�ǒC�&M���L{�����-��	�z �bS�3��g��:>�F���|h����B�|�	Nn<�%]�b��;�t�Ӓ{�����`<�\���U�YP`�2������e_�w��&��.����&j4k�w�e���kQ���CH-��bi��]�d���ף%R`ڲh˫N=~,7�k�&�����'K�l�S�:o�Bʵ�5�Uw>�2wԘ�7���� ��c�ۥ5�~i;�?���6�����u���s�!��,&`��<#����7qRKa��ë};~�n}��(���J+�	9^�Y-���e񸮯*~�.���i*��k�=,˾@j^g��+�=S��sX_����P���0N4�� v�x�ss���.��O��l��x�e���8z���(!I&����L�7���$:^��^dN�-c�>_�*�������Y�	��H���H�	��e��x��@|�Ǆ ��4��u��::%h���b��A8�|��R8�r���l[z�+	�n�x����,���|`���]�f=�\E��c� 4�_�I��a��%��nѝ��p� "�-�%E������1��=gbW� ��$��vW�eN(l�"]�w�ivn����+��������U�r�����"�趕M�H�\ܵ7�)z�Hp:M��	7*Q�p}"���҅E��'�[u�o���3��VZN��.֢��KZz�i�ʝZ}��h0Xt���~H3Uw���������d�o>�e�(67�W���k��rºU
}��jl�E���HͰ�Ҙ�6�'%
}A�poU�#B&l]'���Ԅ@���*´���+-äH?V�}<e�9�κ��gi�4�b����N.�R�Atm�3��C%]����Kh}ՠjȱN��~I��,L����tN�XO��?�FYd���o.ǲ��lX+�<Z���?�ДZ�CSU�8:���E��8?'�;�4��U3Z��,�����_Dn��������a.̂]�t+�,ď�������<�Øe�t��𮫝�)�uL�$`%8\&=�飾�S%�	�I3��)�m���m�l���}���t�Þ���D�,�,��i�C@x"�s�Ϥ�ݩo/�D�o��h���u�e��P�lX]��Y(��#l���~f6w|�v�FA;y������`ל,ׂ�4Gh2��SPv��tܓ�>����̣Us�~}�#�A�0Kg��F�$�W-C�N�(�5�5��}g���Q u#I*�-��T���T���~�*{ɼ�;�h����e���!��n�#y�غl�^��hQ-x�'H��p+��}C�[H9��2�/'^k��~y4\[��R���>i2��� �xږ�Q|߆�n	�o�ħ�L���^�b`_�<��=_� �����li��O[��Z�G,�1�G���~]�.'/�"��	�͖$�NK�js�>�{:���<b�'ԭ�`��z��#���`Ț6q�=������4U��[��
��)\�X�@������|�����_��d��\Qr��T(&8X��6��@�n*W���
ϓ�Y��U.�cܸ3d�.�lqN,����<g ��.�����ݞ�N��&-��F��H�\��#�̧������J��-=�7��s���q�2"<p@k�1���S\i��<[}P�r?��闌IŞ����!s�g�3*͜�Ʉ5�wp�5�A��W��c(����W��) �R텝�yI%���蓑��[;>�8�BJTLZ��5�(�#-�*z��y�	�D%D�S�>%��*�gk��Z�d��|��$�Z�t����%^���1 ��oWJ��W�)���t��t������f"�ҥ3u��vܰ\��P
%e�A�&�,��z5ҵ$��@���f8�ϓ�n����/����D�l;��'l�,K�n�¬^'r���_Y��(�J������V�c� �q��Mn�8yiKӞ�%?꤃[Ut��(���%{r���«�7ҵ�K�gмh�{y2�k�.M��~ؠǤ�)H���恲�	�3qP�n��y�u�
ے�$鍠�H�D��"U*����2P���yW<O���D�q�+���Z"J�V�������Nl��Q�Fb>�R�[B��G�\��`����PF�Ձi�wT�ПS��a�DC�$�Y��K�Ts��	ՠ!�S�YK��:�wn�_�o���"4��Q�̴-rα���|��͢= �J(�e�.�^(��ۗ�	"��`�h8�X��ҚW���R�u�"[H�Z���L�d�R	�<6�%��̴e��=������X���q����9�"1��fF�j�P��m�λ�3r�[�W�(rB��dJN�K�o�ֱ�FV9\��|�E��*�t��>���ĭ�']0@�
������o�N�K#2$U�vR0�A�4z9\^��yr]�-T,~'�Y�t���pr#�� ���C�?�?��Լg ��0!�����5	ʛ�gz]�g��%X�Y|��2T���du�zLz|��x��KI���3u�Mf����kh���!������n1��ڞ֒WY��4�I ��ԒM��.Th�V9�̂���kd��E�i�᳦�R�W����ἑMWP�v�*�p/ �gmɥ+�S��=Y��O��=ԸW��dM���{�`��7�+��/u���:�y�=��DQd[�9O��
�g�sL�� �[E��2���&���ю([5m�ȴC��#OЩt�2��R"�;�blD������p�}�4��]6���yie}'cD��y?86��USZ��1�쓤������{u�����ͥ��=��,�p4?��,jD]#�
eI12����� �d�}V�L�V8����MA�pB��+�1�Ν����|M`L|{MW�?.�RI6j�'���81tM�а�Q�n�Ņ6��jUS�%C�6�=�YX��ӤJ�(2&W��#���#,U�� �)��;?[�]WpQ1_��Tr�-}�x�d#��"�뼿�G�W�Ƚ�A�LL�[
�R�&�X�En��ޅ�]h}���ɢPa	lI�]dۺ帵$�z���[�ҩU��׬6G��W�GIN�������W���'���9n[����b�b���g1,:�FCL
��Ƨ�@xMj�d.عt�A�Ç��Y,��e큡�\��ir4q�"c}�r&2��*�Y�~��f�ir˝JԞ�v�W!���9�,����SL�zr�q��{�~1YNE�����Z]񫥣���K�j% �[�uaFP9]AV�������4Ε`|3�j1$���NqӴ^��^��8P0��z��{*�?|�:U����+���{P�0���
ߝ�d	1�60L�q?ꊷ�mUP�=);A�d;c�@؀u�눚oF۫�v*�!��&=�l��d��d��d=�����������[�\��L�5Cc�9���R�� \6�@X�]R�Y��_q��reDbs��C�T�-��a��� 
"#�PyȰa��K�W�:Mk��
Ĭ���dІzA�Ԓ�>#С�� ��%���%W�x"i^����8�=W�+V�	<��cP���N�ͨ���O�>%_�K(*XG3�������㩖I����己�^t������4d��!��oZi��Xχd�����O�Cz*쩤L���W�Rk����u4d�t��s�D���%c�B=Xv-�z���Yɺ�{2����TdU���3����B�=?�e�실я�V��:�_Im�@�T}�~-G�[F��[�kG�s]�$���	�]U���M�f�v�0�y��78�U�w� ƸGQ�y���N���ߋΩ��&�����k-��R�;hI]ĕq�� F��BU۵�D�b��Y�u�����r3�Qf̜/��;��e�G�4:\=\�I�Y-Y-("p�/P�������T4�`����@�K�!8b�ү�h���>���J5Fl���ӹ��8ݬ٭�I�	ນ%	�����y v�����i������76��酷��2��o�֒��w���;4�ڸe�����VO KL�@Rw3��=c�d+XIȮ���2�n��vQ0/��`7���%<���35������7_�cc��9��r���n�o��:2$]; �79��.V$A<Q�G������d��_���x�C������zZ���h ���=�k�U��=����	���8AA���Jس����,wO��r�6���qF�hᴰ�C�1��8m�Gy��L+A���P�\����,5���㛵��z�8p 3������d�o7]�7�la?��0��w�t�?{��lv�O��kd��so�rm/��:�J&��o5e�T�g�iGe��/�+�ɈSe{�)���ن|.�ӳ�!5X�ӵ��Ag��|���@+����Y���"������)�=�py2�������/�?L��<�M����{F7���;���x�x
�H.}�*���K(����"H����{�'Ұ_�B��ml@��D��о��&�a�-�K~S������t�ͻs�����N���R����	�����Ѻ-��"�� >��#x�4��GY�Z�ӹ���j̫�[�W����qE`����U�Q��}/����bM��|���Z{La|�Pw�ūmgaI�w��x;-&�M����jUe����;��T~�ۉ���-h�ҟD6���M�$�{�]����+����Y[.�M�G�Q���*�˾��݃H�Y-��.�2�"Jx�Q\q���E�8A�)|�i=aeeM��[t�Z�Uz�����x+Q�TD �O��f�蒫�[]�&��~�XS���`�I�Et��+AplЧ�$����h�q�[�W�&�#�:)�_$���b���9>y��֕���XKY��ʥ�GdpX:�V�]N~6�Y���k�e�ǟ�Ȟ�5|I+&���w�ٔ6zy�,(2���skkB�h�!�Au�.iUh�v��k�}��dA��J�����Ă<_���45�iQ�6L�5�~�շ�:y��T*v����@�Ko���.\f8�5΅�!gX�R�&ϙ�_6d�3{�*�tfh."U,���-'�ho�Ӑ���D(�8�H��������_d��A�(�x|jU�zO���7'��$P����JG�Ajܥ�%���:3�a}�eS濽�[u�G<}n_]��6#�cp���KT���������nN5�i�>=�����WcQ��R"z#��#l�����ʾ�U�$X>Y0CM�w�6'�` �7�q��i��<��d�f��aS�s�:���'�ZPG��<���~�Q�&������O�lcО��3i�5�#��$N&�YC���
��@��g�$�J#p������/7Q%���)K����O
չ��k3�"W��c�-bQ+�����{��Ґ敢�Ց�|��J�;����A��#�g��g��^� ��9��l�-�ԇ� ��eV �o�.�{hl,"���?/�A������3�J��X�$������!�PܩZ��H�-�%�udIq�[�M]!�eP1�D�z\c�W5F�.F�V��0�\�i����1i�!�{Y���AQ�إ$��ô*��S��lH萢�vA�C1��VX��,c��3zM����:Jn��4�~kB~fʴ�r
�����Vj�V#s���J'�#�p�p�[��50>>���R�.�'��ڗT�V�����!s�g����~���"5��*��0b:�	�&�3��u�4�r̫i}��Uhփ|\F�%������ Q�D@k���ܜ�I6��#��ю�4'e���K�ÕH��؎�|�4�	]a:t������Z|#"�V.�|k�2�A��<�O��'VL?b�;g�Ͻ�s���̦L�(��T0W+x&& qܞO$�L��6:}i��U�&9b����k����oƥ@"�O�@����1�"=ו�
0łt"|�4!��!��Ojk��,|�X�ҡ�����)���~֫����g����$�X_$45���3������Zw`i�����@�,e�՝��]$^!?$$mMц(hIi��������1�����;�ō��ikFH��۫�y��Gr��bp�ov��tEǣ���w٦�qI�1��:�F�h
(t.x�~�h8�����2�w|��� �9�Q��R�|K��^�"���h��2ۯ���649+KC�Y��F�I�����n4��Ôڼ*� d��T�\��˩A�H�9Fûzj�,N
�n|%AM;�/�`w�':Y�e[�
(Eq~�� �a��]��v�{���oU��`!��8y�%�J�m �����+XlxVHYEB    f314    1b50H��4�B�%��A�nX��IX)�pM�������%��O�Ǽ��I�F�*��d�%�@�F��TTO�mQVb*�͝�Ƿ#��'6��&�@~_Y�>�#|b�(�f����eryU�0<���O�����L��b	r��ZV��d���=S�6q�o�Sq�Ó|[�@�߲���P�`F|��z�h3��w)/}n����d�O�k��%���5B9�����*{ᛛ�%)�J�Gb��no��UW^
u��1�.�"��~�=�A�'9�����P>]]����^g+T&J�.\�+J7b
�@w��Iv�E�p�~$��|Q�	Ȝ���XB�0�d�.O!9���9��;�������MFe�N���)��d�vg̛��\�Q��MA}�&� ��T&�b�t��5�a���U���b���mP�:fn����۵����c��*���l�j�׿)H5�L��<����{� X�\���fʤ����&C���1P����}��_�T0)�g�&t�,EAC������q�h�"]ȻX���_��*�Nl3��(Ľ�O"]H[ȡ��"]�G��01O�86D,���*���|y�$��[��HH�ʨ��o����Ӛj�����Yc ��k�*�K��Nsy�
�2+��U���yN��@� �aU�c:�G��J�$|�_�*�>���&p�H}��u�S�rj:]>��兩I`��-�0n�N1���;E$X���Npe��/ OR���eJ�����8���z��k���QD���Ro���~S�l�s��ҹ���|���g�%�뛵���l��HBka\&S�hCD	+�[35U��SV�J��b�ѿ���e)D~3!����a^0����5�W��Zȑm���Do�% ����N�ee��7��o�B�V �S�-4a��c�xDP�Ɲi��hHL�x�|� h���V<����7���ErP��Ʈ���X?�s�z�ʭl��sۅXlNz�X:��꤆�7^��;F-Ђ��R���RȁXm!%�0�����uhr��t��%Pz�I���%l�m�	�С�l>̺X����4�*t줤|���˃j��\2ȴ�#�}bfv���yKz{�Ȑ���b#�ylgx<�ϩ���n~h�}�������Ў/�|=���Z��O#�N,�]��FLH��j���C_UA�>��隱 ~�D@���h��INUrf56����v����G�4��9_��;�fC���pi;U��F������ պ�}����`i�>t2P�Sn�6:�@i҃����Ӥ��q�py��������gB���8VՀ#?��s�j��71:u6������@#[�����Fs�P\|ˤ���zu ����(��WC�$��8���*�a���(HW�;w��~�l�h)���'��;_��Qf���_�&#sb$C����q@șL����Z��2J�[
7(�-������
��ҼD���ˣ���}��!� *;� Y4����61�O���\L?Y �MdɇP~d��sޙmb�x��V�+=;߻W(>DO�O�� kX�$��U
�}�3%x?��m�h�@O���ck�.��mPI�t[g�9��^�!�}r�!5��B�I�����+C}\D��� ���B�.ѵ���ࣷ�R�@����B4d�HnП��E��9�BK�wi��|����;V���4E��/�,���"�6�0�ǹ"��4��٩0�����G������V("����k�BC
0P��ƒ�����H,�?�����P��� ����"_X�󏦊�z���"ފ���X?k0�`䣋�$�X3tA ��bS��l��Gk��+��Z�%���Z�,U}n��-1�E�i3��Љ &�7ؓ��Z�uk���*qk�{����ذ�&z�d(Se��!�Foi�Ѝ
�\�~h�K�r�q&	�sn�e�U��s�����h�kY^�u�ǲ�,e�����e��`�/)���q.�c��Gjl�m����*�5�lhTa��3�qXNrbr2�R�t��-�eP)��Jo�_���N�go������\GW��U��u����[CP��UkvaϩÁ�zX-4��$�yK[ vO䦭MM�����z��6t���ǘ�],������N;_��j�9�P!Ln���ޕ����*7�;�{��165��כ��!�)Q�@�`"�Z���X�q��i>t�,\�@i륱���`?6X�Ҏ����no_����tT���1�\m$CP7l�w)�6u�@`��:U�&�c�^8}kL�c�'�d���(7ouQE�[�̒�r0�3����Hv] Io�m0�Z��(�q�g�0����C�07M��)���4��9�^��5�
�؄s��-�?��./X&BQ��+�+{���3򭽒�4�<�0��W#o�Aٮ�y�l�� �.��ʻ��ipMl��kzݽ+��̢W̔B*<�.�i��@=K�6�lI�z��ʱ#�_
2�Aj��%��/t�*r	v%���f�J�!V0��ޜ��~G4+d7��M�W`v�yK;	uH|1dل�xT�C������	.���dr�O#<��N�[�~�K+
kM��`�ܽ��R�u�Ҍ0.��z�{�b1�����oDY��Nx[�-@�����K�V��U&��swy�d׃O���pY�碑�/�M�~cTOzZ�N}�H��'I�#�],��UЌ�G����4�3�V��jY;I�1w��gJ⫥����'�):NQ8�������5Qs��ߌ0ɻ�Q�UD��1�P����A�,%�e�+OD�w�éę�Ҧ�:ΗuÁi��j�le�~T� �`4���mN�E�'�8(?�ɵR����ST�;x
(G|���^hiz�:��/���J�n=6�?��@-�Y��$��7յ�"v������x��<�XB&h��R���^?EE�is1xsP%�&�Q7Ҹ1з2�ԩ-sƞ����pЮ����������k�1�HrjH|�d9R.�l;��2ї�˿��j�~��K�j�>�|� ا'AŉL1}g��U�H1���pw.����2��Wq���|*71���v���	�Y�
#�R�g{�� �̂��G����׿�\8�Ԭ������2a��"�$v���H0���#�?����&��� 7�7P_�Rh��h@�1�Y�u7�������k�i�ݒ����Yd)J:~YN��Q��
e93`-Z��s�B�����ӂ̆��<*cK��5�Ț�e=X��2�5e[�1d�!��=A�1��<I"\
<��X@g{]�u�p���T�rU��]��v�	~"bQ)U�����W��{�|���F�^����M�,���Q�K���K ��b��r�&�����Jc��q��O{-�m�p?����-��½^T���O6Â����U'~�/�XXT��;v���Q�7�k9���5�b[1�JUw+fΠ�׷��>����$DQE��b����?I�"��tO���I���[d��)��s�ɐ�DO��	����lG�yNB�.��tJ�;W'Λ��8�+�&�����-6��n7�)29ch֖v^����WV���a������3�w�d*�ܧ�L���ې~cG�������Cb|��:�^��}I��/n��q��S�+�h�z��9����~$�о�<�-���М�$���$-Y����`?���^���(n��[Sc�1�[K�d1���?�H�[3疓�s��+U]��y_�*4/ݷ`PT���^�nQ\|�R�P�H����
粐���0��(�J�6�]ױ*i�؃�E��jL�*�]�\�4�8��~���v�ˍ�FĴz~�&��!�s9�"ϳ�VƱsѪQw�Qj����јZ�a;�mS>�;��Ep�3|���8��wg�ɮ�[��Ydo#���Ll��z�V5y��s�M����A���& 0��%[ۼ5��OZ�e�$@f[�%2U�L�[n���F+<���1��Q����zH�
J�3�gR���$�UNI����I�����QM��s�e:N��U����!b�qб1�������^��YI3|<��͊^�5)�[�z�&��9~s6��͜�~�A����n�1 �|�%����!ҥ��0�/��5��f�'�ڄ�d���n�{�}����=�A,bO����Fl�����)@U$(�(N�P0�mmzЯ�:��Ua�
d�v'\Z�:���zD����������<��c�[��=�L�)[*�_�"HG��H�<��z`�����4��[1�*�W�ڠ�*�v+A����7��S�Yw����{��*��I3T�n	�@w���r% �)�H ��]�>�ճ熱���ʪ'nM��e�AN8����ڼӘ�C'�DoҸ0q���J��� 0������<$	���{�h��n)�Q�`���rva��һ9� �}=J?a�Hx��#�	��}���o�.l7n��������-��ɤ�ޔV ��;ǡ(�a���5�n����yt�����J��0I��0�BD�dݜ�f�e�o�4��~["m�ej1�ơ�{FZ	�d[\H�?t0����E�|=�UAa��|$*;;�'_o�����'��<G8BE��#H��ƃ��gWl�9�
Z4�v�P� �P��Fw�ⓋU!���>�/VU^z�����n��A(&��܆�$+�a2MXa���U�y�(��?���WO�3�,P��u�$��'�u+�|E�:8>�7�`U����ؔ��F��#�M�Ye�V�H9�צ�_�pS$��{?x�.t(�Ŷ�iI1��P`��г<N�lp��Y#�)j��W3pg�F=9�����S"���u��9xe�ƾ��V}��]�v�k�-n��V��,��"�3m�\�x�ނ?I2A��>�c($�j|���|�����5�u�B낃��5g/ϛ����8���M�m�n�����_`��o!�q�+���}�*��no��Z�c8ZAU��}�a�-yY,�YF�@%E��[��P&����3�ﾝB7į��3�h�u�ґ ��._|��1�햅DAb����>��=��%�c��G(��}���&��.�l��9��-D��0�O�(�)Y>slI��9�3�"��ӕ@��ކLn-�j�rRq�����pQ�I}*>h=�b�Y�L}ۋu��Չ�Pc�!�>�rkh��-�n�^ �A��c�ɨ|�Ԩ��D-�k�&{)~g����X(��;�,��b+`���W��c���m�!�jVRgٜ�^��b��NE�T�J�b���W$�H�[�󗮞��� ]	<���bC�Py1'5"�M84����
Fi�3SS���i�J^Z��Mdե�轏t͐���:���S��G,.}�^� I��g;��E�z4g5m�l�<��5�C�z�VZaόv~Gym����>oV@��� ���8%Y��o��1p��=��Eb�������ީ�p�Z��~(��1��T�,FyrG�:���-�`D�:�Y���b���d��g#�����/��� ��ta,A�K�*��k��g���9`& c4���cs�h�����u^a�l=��Qd���E!��"�5��#�����R�G��k�j*BV���ku���a����AS�\�pؐ�:�`�kI9�l�r�z�WA���T��/���^���:ŸZ�f^�Ouk���϶��,VX�2Á*DI ����B�!֯�f�{������d��\f/�<�Z�F��j�3��T�M�jLt=R�Hp�$�>�j�㦐E�8�;��\D�� �g�ͤ���@����yҁN�^o�C}���`��3�f���2X�&�x-�猾&�ש�ĪX��z�
�CwB��g�6�V�q�|�]Iު3�Aն�u�r���53%�i��mW���=���+�������-�.ds�i��!?z���t��H�.
^��-N*�Z�f�Oe \�};Rh�!��y�2z�@�f	E%a���XF�N0����5s@Թ�Z؃���Եm���j����ə��ֺ:;h����=fiG���D)���rz�#�qN���Ĭ|L L\MEK*9�ǱB,�t�k����_ZQ#��*o�TCQ �u�h�����D���a5+gP��
2O���Qo�>d)4����6�)�K��8IP�XĆkKw�k�p�*�΅r�m��S��UN�s0;�U�ߒ��R��>O�,�DV�"�]2�L9���DBs����rr��Y^�΄��/�;�n�9$?�X��p�\�Õ�8cn��N{%'� �&1\"+Ba�)+}�P<�b���ˣ~�������\V׵[�eܸ�P�?�X`�N����Q6LA�4_�<�0.G��,��oӿRw�b����a!��F���$>bX#XN���媔�l�U�s�I�h�:�G����7�BY���,zwE��H��&&R�bf�͔�e~d���o[�M�IM�W�QK�W
8CP9[l��a����%΢�	�k�u,V&a��{2��}�,��VL|uH��
�$��bAG֙^�xSA]�r�V<��j���@�˷�4;
�ks���+M�gj+F#�)d�)�î��"�W���3�6W�%��h�:u�r6�l�V�&xwc��A�\�(��Xi��U�2�� x��w! G�"-���X	��n)��/;&N�s�5g|���^����^Z*��]�зEf��B�	7��Β��B���:��z���!];�������{ׇ��_�{(:X��P<+Ȩ��6��lsTQ�Al�D�e��Vwi�]6<&��H�ؚRo?}+]��E����}l�GO�