XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��yO�T�-cx��K&dޛ]��,�R$[|��	����5Z&�8��9x���0����aw��lI��)����ֽ��D��}-�G�?�l�xS L���p�79�xpF�i���n^�aO���YZ���Ɍ�Bk�F�]T;�k�l*�����7XyH�����=&�������wi�`���^)3jp��^��N-��׏pB�l�*A�.�*ᄆ|�swOޥ��fU7���u��b��a������A��k�Q{��l��4�����c�o3���vI�SZg�� K��v��6[�ӎ +gC���S�#�M��!7��Y���g2
���C����Mؓr�_�m�<��5����o�K��|#?�i���{�Ql0E:t��Q��7&n�LЀMR@�h�*��Vt�~͐C�����
�t��w�i�����r:�B}wX!TlZqxGUҿ�W��}$����2Y�b{'{tX
�_���XJ�򦖼���M~�7!�'ʬ�\��>��U'Q3Ƴ�&� w/�,�6�[�U�ڸ�ns��"�.$䢓o���)�y;��ezi��X0����/�.�5��a�ލ��4K F�:���m��n7����65_�Ms�����f���:��o�����e�Յ�.��p��3�E���ڜ�m)��"kl�FCvM": ��&�$?��Ô��4���gRX�$���
�μ�~S���ri)�y�1A�\�Ã����3LH�f:*��7=��^�5v�,���G�r���5��XlxVHYEB    545d    11d0�ː6����S���9����^V��e?�-%�5�C����
�J#����9�W��t������Xt%��^�1P3��7G)f[������٢y�GXC��/�Q�isى@r�����Kh��I�E���L�F,4� ]��ߛ̟E_C-^mG͸ulL25�n���î��Q6?ot�n��y�7U�M�f�4x]i{0O��:Ի`�����6�s�(-?m��&>z��Q�\-P���4R���v��h�Gۑ:�-�s.F�Jd�$�+�/8�k
C\$
袤��������kT0�����#T�̽�|J�%Y�d�52��]w��Y�$�)E�V�E��u�+WB� ւ�x����� `���.�͞���2�k�{����½*�Q� !�+��옟;�ws�_�2/ο�6�K�l�U���
��h���������Di_��6���"(�MZot�}�<�!1E����!MfF��M�xݮ�p�M`2���_�r���vϳ:9�.�7�]�U=�1��)f�	i�:�_��0Im��6������)3�|V���l&���WԆ����>���C�x3.�����UX~!k������e�� �֟%����ξ�'�=DkslM^�"�	X���$�_"wg(�ӵՉө6���U�'������Șƣw���}<��&�#Js"�&v2��2p�]�ר�J�g��|��᛬1��j�&P ���Ĥ_��`i^6lS�B/�����0����+����a�)׈u��_.�\8!@�<'Ӧ����E}Ú�rZ�gc�4N���`Y��n1� *=}W��� �{��a����B�}nJq�j�BNjo2\�ڪbT�C��*/���{��Uf�Sh��7��l�y,��G1��X!%z�f�@�b㮜|Q�8&��P�^]�ͺ��d��]���_��C!h��Eb�g����C����a��e^�����y��41�|KvSZ���@a�:��(�(�5���5Z�$�����Ρ�D9��ZR�g��������y���ZD/$����a:o�x�% ��/a�d����:%�"�+�[����i���0+���<�PTM}�,U����U�x�&�?���*�ϑ�}�A�^Z�_����b]LI��4W#Z��LҌ�#7Ɂ�J���g"�R�6i\)����y�,��ͭ�_,������!����|�����Ln���&MoƵ�`[��߫�}��4��R��;��۲�������0U�n,!�/I��<j��t߭�Z���g ��b�!�=l�:�65&����6!Y�2oW��d�ܠ���'�0؇��	}"W�;mPGdNBE}B�j2 ���֞��E�'�e�������K��@�C������#%�%�O�=��
	LB]���l�3����� ��S��9V(�np�k߼`d���I��NxGy��C��e��j�O�t�F�F� �`�W�#��[csЧR�U�#H�@�=��:Z�|�<�#�u�p~+�Rּ���u��8��c�'�]����`����[�b�䇺$�;��P��MKqk�IN#��J��m�Y\K"��]�&+k�o���Av륱S\��9���>
�zk�>�s1��\��x���y0��nb�7����)w!��/^qGZ�@�F�fGp�)FJ��-P���fG{�+�<����������ct��a1�aX��w%u��#�ZE�f���{�&�?�8�Fe@������A�%.6,���d08�����<��
��W�p'���|{�qdR�ߏ������\�#[�% A����$�}�hkR�bL���-�P�2��LW)h���]��l�{�374}�%��}�+9�y�A@���]��x�<y\�t��������4��{�7�D/]a�H=U�S��ũu�Vؚ�m,HP�*c�M^�L��`��	��ϲc����7iAx%��o�*�b	���KK@�6���T�}>�v^Hr�NT�$	I8�g���.M��:�W�n��`IU?�ȩU��,��D���2�A�U�~�8-�(F�}�?؇��7���c���>�2��e1zU3?�i�{4�7�>Ry	3K��;�_�N���|>Xi�=YcWU��
jMh�x�Ҷ��3D��ն\V��-�y��ImP�x�yؔ�}G]�Z6c�X��W�I�ouT�F �[���\5),9^����[5�qv�#�[c�u+S�(�^��N�>�8�v�u�Y�~���)�J�*��uADY[#�J�*L��'P`8��C�&x�2{/Ph���n�
��r�����DξHc���:�͗	�&�U��-���� ����[3�u�B
6�Ȑ;�:,=<^�BY,��iλr�Z�y�+}�=7�'�+y]IJ?$\
��z�ʭ�Y#�1B3��re�I�%�s�Fu�����!-��C{($>9i6��4,���5��a��
%���
����� %��v�q�+��P�p����Zb�j�f�g��оެnL�VJ!YU΅��e&Ye����hm���6�$.��0ᐅ[pqtZ"��4�F�|%�r1t�0��c�� ���5v����8����B����`[O��co�V������i·%��_��]
$���<���5���w��4�8-&��!�p)�^rA(Gߍ��|�h���Ta?0�~4�9�]^ݴ~��b}C\��PQv�$�gM��b#72�X��}������ʞhhM�T�����ķ-Yӡ�`��Т�_��P%DS�F��ȞtL8�?�^8���Ǥ��$RWCο������%p�5<��M�
����a�\�%U�'��\so ���U��\v�tP�6���p�0s�8�^���Ӑ�
Й�a�cN�Q
7:�Ў����[����Q������,vC��?cO�bL;�*�v#��S�(�gQ	�2���+i��4����B
��ŞD�{/k��4Fl�kT��"8����%�71�%#�Z��X����y&8%�e1�&���-�~ͫ�f����B�ef���3���2]2�օuq���өo,���%
�/o�S���)R�1�iʲ���,�	���Y7+�7?.W�8�xٺ��V�m>�q&�`/� ��7��wV:� ���r=]AuP��Z������3=Q���q����-{�u����=^�TkvZC�b���=Σl
����b�-\���=3��!�s�p�I��>DYݿR�%hX0Z�[�n\�\�AF�:.bk�������:��=�?0�g���(1+	WoxrGx��b�@t���_�����������6U��Q�*�e�qN���2�����45�o�^КB�6C4^ ���� r��)2n��Z�R���}�Hʙh'�����.z�;���dx����s�!;��)��g�3Ά��x�F�+��q��@q������ܸ�>9u� VԊ!�)��	�x��y��zh%w1���1ⳙ8�z�ܔ�5��E�ȭ):Ѵ؇��i�%E���m $I��͑-		�)�}7�p��1�R�������W�Y�ټDJҹ��#�^�������Y�7`���NP�yOO�^����S�k�M<�Rp>@��xb�J*TC7��b��l�s������'� ��C����� �*�\n�s�6jC�K7R6��ݥ[L�o�*@e�ؔO��l�nф��϶���Ë!&�Y�B�����km"��q�ĦD2Z�h��WhM�׉Ȣdg:�&G��"�_�(��������,�9Ta�!�9�Y���Xt��%$�,?{/�?I��2������LO8���V�
�����P��/37�$��nS��و���~yN�-�/���eJ�E=Y�N���ƈ�+��?'�ta������Om��
Te��r�[�^B/�1{�V��_߸Tt:$a�ld��i��]|��[��8G�=Q��;PAB�
4kƺ�c��$��|X�',KrO����t��F���4�h���a��7�
���L����g	�O�>����dp���(>1���S�qf�v �P)���&�,4 �����E^a{���(�˃��K<��-"s�$�V�ĽS��G~�,����Ԭ��R
#�Q=@��b0|����
�;�nJ��"xQ���?������th �M:�ϒ��@9"�����>���ӯ��v�Qc$/H�0��4�ϛq��� 2M�:�Fy����'+�˛�V��T ��B
s <Q��d�(b1��.�&~�r�E��U"~}W�6�ST���t��9nL#��َ.Ω�O�kK�֐�)�U{�:݅�����������7%��=d�2�iA���Ãc�Av̺��Q����2�*�5��S���aa&Qo&���y.��D>[�y������Ecg�i�������<a��SP��hJ�"��oޭ��
��L�on����,���E�}�)�Eq5ъ��R�*��y�	�>P��m�(