XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Q��E�X-	�PϽ�+����:���^��)i�{��p�@��b���~, 0��9*~@[�{��ENhe�pW�M���T:H�T����;����S����3���I��iC��\�9ɦ��}�ǖ����eK"(�+&݇�g��O���H ;��~|e�:p9��^NZ�a+��$��nw�8<šV�I��������%J�0�N�ӝ�Oc-�lO�y��lW@Y}M���`42�����E�s${U�alW����#�R�;\���t��q���4�zx4���qIR^�����>oM[���_|ֽ�8м�RИmI�S�%qM��p��/�����fuDGR������/ �n�)�d<���{ïN�Y7�RK�7]�^_a�hU��#s��4ٙ���*�y�[Um������˒����� /g%? wa��B����S��4��ng�d��[�hi��������C2g3'��P[��j��.�A��Z~�!�����������0�_B^�ƀH��
��%����{���2u�b�3�P;����8�C�S�4tI�h�oxpf���)��n�sY��ѽ�Ͽo�t��t%�ܱ��q@�4�\3V�8��Z*[{sKm&Sr�3�aB�m9���S;g�7җ��x�8:]���(\9���=��>yw������r�π�ҷg�(��/TH%X-p!7���z�A�fOb������*�����#y'���Kl�o=+�<����:�2�B/3u����, CXlxVHYEB    fa00    1950*�<��-���۰-���p�&l4"6������c*ō6��]h+�����;ퟝ �yU�ۗ����@7����:��_����7�~��8��LXa��dp�OO.�|"7�[Y
Z&���h)��݉JƳZ�"��gaw�a�^�r��0�S�y�Y�G���=�I��ބ���wh��$�mj�A�/Fk�j=���M�7�(���m�oi8�ZW���5j7�\֮f)a��6�唪�0�����h���#y��<��@�n���hl䝦��炩	��͏;�)~3 ����#�������s�Ȑ��L�1�¥n�:Į���2�4H�P�$E�n@k���H&�:k�����IF7�\��oTS�������U����x�P?�7�	cLo�Y�͟l�!
R�G'a�q��"s���e���K��X��#�Z�=t��B������D^�{j����r��xe|�5bm3��4�����s��f��D W��DK�<��{Sgݯ�YsD�6���AX�����'c��Gj=�PH\���E4aY@��-;�V���:\�D�/�ٓ�T�.��+��a�C�����M� !�m(��rU:kۃQBz���iU��;�������}��	�B��@�'Ԏ��(�i�n��p�q�������OyF�^���ֈ#�PY�PH�t�CS�e�כ�dǾn���Ĳ��`a]6_H�YN��[�u_}UU`dG���+ɭi�7'�3�f<j�G�������ޠ�G����� ������g�{�jiZ;b�N#��0� P�_G��¯Q6E��X�8Rt,9�ƫ�t����C�o�7od��	�6"6!}Lr�>�~�~y�j���<b����2j��~l&�aq��(@�N%k�藑J����M�Z��~����c��'�R���<�!�q��C����E�.p���z{:��S��f+}����
��i��C&�Ʈ������"ղq�|�(T��!�2���4�ȴC��jyc�l{�ݔ�vy@������k��u<�R2U�F��q�j��c��!ep�j�\"d�]�
��c)�����E�C��B.6N��\��ʷD&�P/�~7��j���K�������1�e�7�OC�ܞ,'��;�����Ք�نLW��z�ȹ���գ=V���f�4[)p7��n�zP��c�I���:nCUU��.��j���:�=/w6?�Ù��(v�l����O�0ݏU{��;fFQ�B\�>�&hr���=��
���U��^�>8j�� �;�P�\����5��$�Y��{������i3珿��������}�G���~�R��"�LR3;�~L�kG�*)�b ���{�����<��J�X�־q�sfU��:�@yp�ggN:�=��_̒�I�p�h�C������v����5|#�N�b��%�E?#�R�$a�8�";�;?��s�+�<8`V! 5�e(X������Kб��aln0hÔ�?�34���{��=iaʀ�q	_i�Y8��	p�|>E���k~H�Tœt$2n�M��;�?�ew dB�f�Q�]hYF���Uc��EE����e�X�r��~��N\�m���[��0-��s�����g���l�Xa�+&U��R��Zr[G�:��=D<���� ���<h"�<�חq�5�]�G�b�왰?oⱑ����쉇D��_P#����H�,�}���O�eD2=�(���N�.�Lr�jzh{���1},�K����X�+�~�����$�vr͍(�%�h�t��NW�o��F|�[�|�a�t��c#6�e��)�F�h��)�~$֢�l��6�K�H�1�� �D�6~����LGa&��'����C����Ƙ��u�i��Z����s�M�W5P���W�� ���Wg���)���,�"1EU�#�ݵ��ݜ����!s>?,�I�\��ޙ����u?y2�mVS�C�Hf�O��T��,v�!OtȪI�Z��ϑO�d�O����m	�;����5l��&|������R�Vb��n�j<H-��hs,?��l�g(u�F:T�7�t���1$��ܘ���h������g_�Vf�S��l��ף�~��b��(Ѥ-����IU�u`�TFJ�bڿ>��/f*��)Lew���)˂X���fEpu�a^̥V��m|�s���^���;`�eQ�.�}@Ðˊu��d�B(X�Z��֝�N'$�؛s�]]!kZ#Nl�M4Q饫>�\��.���L�u�I�+Ij:*��(��T�����G��)r�mi�����w�H����ڨS���.����6�������;,�Bb�B��Bn�IEfL�Y�7��N�)~ tw��i
��Mȑ��N��b�$A���4�����"s�_��ܫwK dw-@� �dCC�,1�� ;���9�T�A�铮\��. Q+��h6�@��,7T��f����8De�x(�
�)��w>�����~�bj�i�w-w�J��g~��յ "
�@4g�J���h�)[J�i�?����gB܍c�Z���.kT�>	SXX|��2*;�)cdʛnLzd�r2Z���3�;>Xa���k"�͡��D����Y�Ol� ,Nh���A����3���ڥ�A�R#�mvE|�;Ɯ�="@�w�@�/=$i���0
v���b��m��ݏ#���,�x-�:�<q���/g�4+����}z���t�ۙҩ$3uz��D*�d�g��M�G����ޗv{>Ye���'kغ���(�+TR��F����`bAdd
�Nb����Հ�i!��񊈉�6�U׿Ҧ�@�?!s ���1-���S"2�bM I��i	���'�b?O�	M=T'P��5?P--��v�Q7�j �����-�Vr�ľ{A�+�6�|���9R�����p�\a��D��c	���:�b�;��>c��G��Δ'�dQ�`T��ϐ�Á�q��i�:�'O��(W.�f��5{{~*.��M��B��j@M�E���,�3�r�n@��H���-�����Vj+�����E�(_Vz�>})�j�Z�D���E��>�{wlO�w���- ��I��ޘSr�@QܳJ�?&l�P0�0�VuY�d�|��V�_�9����%^����]q��o�W�*\�����"H5�J��LH�+������l�^�=>�6�����3#ǳ��s��dx��G/�'�\V'oE\V�MYb�,mb��qR����o�������隆#��
��yi�"��IQ'r�Vuw�&�x����Fx=Rq�q�$���}|V~Uʱ�Չ���Б'F�b�ԫ<Z>(\��",qt�L��oU,| �c
�ÉQ����z�]U6\� ���o��rh��N��.hH�	�Iz�4cz�(V���]�|����ߗ�{�%�EiA�^���,C>^$k1g�ΘZO�d_9f5��� �V�L�"��b�#TS���aL����V��L��r�!�G�5�=tdĸ<L뒘[-q��π5z`�e�y��!�w�ʃl$�TI�J�Ĕ��7�`�Y巂*Úp�!	E;��Y�=g��a�4 �S�3��F����hR!c�>'�'v�g��ƯP��L��H�<ß���#���o��Tn�^h+N�<����9��K����<�}�=��M������m�ʄ������>#�}}��Y����N2H�ۋ���:@�|����q�� ���3 f��0�%Z�+�K=�˧���{��s�.�Ù��vu+�6��tp���Z��D�uJ�� U��c��x4���_�,�,3��D+Ĭ�?�u�<��n f]<O'�$�g�(��ør2���;��U>�as#h}�A;'��I��QFY(J]g��zFj� �K��-����T�d��L��� ���b1]��*��쥑��	�a�^=�]����I�<sEM���w'���Nq}� \���'j����c,���Ŝ�#B��b�������\]f��>�t���^>�8a��\R�ħɀ�㨣UJj�1z������*zK���`�?2{��F�ʕ�I���dU��H�_ܓGZ�<�a�m��V�ާ����ƅ�6��/p���ﺎN�Ai�`���+I1�;,�:o^�V�r��׼��C:������!��A�� ���¸ȭʋ?�3�D$9}e&����n�(�t�ıDR`X!ER~�A.������{Pv),��.�`��  {��Md��êU1�E��jME|��
ݬQJ��X�@�.@�?�-��@7��X�@��Avq���=�2�cn�Ϊ��^0k�=<�����"2^�v�tk�0��J�RJ��ev�2:bU���FE�ӕ���!ת+iB�p�JM�
��2�y��3z:K{ ��B�a�����[
u!�;�_s�Z:q���ϙ���ϬB4�{Q�)��R���Z�����X�Jd���89Y6/� s��A�J�I�n�Hk1�W:)]�h�j�{������|�ܢΒ�+E�xks��vC�͸���LM�M��E1�>7����;�RO�Y�V�ZGv�%=�ѺJ,�0�1���eC\۩*>�?��/!�ڄ�W��c�p""�@,� "���a,�y�~!�饹C��lOE/�sp�� Gb�C�]c�掑��ɲn�8s�wt����lc�`��I���">�4���0�/�$5to��Rf�=d��*,���P��,�`Q�Fϖr��S�*&�K�d3��*X���J�E�H��$����<l�\�"Βb��u��ž��]1Kx5 ����ۧ��@�Յ~i�����>��৭r��"��O��t+8g8{9H����>���������.��K�����W_-�$m��LĠ�I��QNq��9����!962hR&gS����F�&���"�
,XK;��
%�"�P�^4���(0�}mos�L��۹�ck%�{�§ǔ}��a?�Z-��7<����*����G:�]��
W�mJ2b�{	�4U�SfCW|���!^��ģ��2�Ȓ޴W�������ïɳ��)>l���0Ԭ�O�zQ�tP��z*>�9D{&���AeOP��>�AOk�gfM��tq���d�{����i�4PTm�,�\��ӏ�5���y��̥z�j���^�G��8������T�)ַN;Q5����;)i�����fc2����&{n��Gk�ɽfD��1rOq�\qo�b%θ���;��C�;����$GV�;�)��/�O�m~����=x8�X�1=۴0�+MQ�O�� bl�!F�c��fx��B�Dok��O����y3�]�={�C�K���2 (K�̣y��U+���6*[" v��L��H��aa8�
�0"~��,��}���!�[X�n$�7ި�-�7<!o�`8�i�xK\3��A5B���jE�?�����&/@߁mõ��X�ʐ�I���K�*�6<
V���fǝ�i���AF��U��t�2{���T���wN�v*��_=f.?1њ5�:Ǳ�<�5O�����g�zf��	�.оo<f%��D9s���";P���O��C2�[��V��5_��èv���O�q���}��?$=z]�R��sOӮ����쇓�l�X�ߖ�C�0}��ܤ��kmaw���7�↔�g�j����{�<��(nMt��[�-5��ޖ�;���4�b	��RA�H�yvѨ�3q��j��M�U֍ĈZ�H �jO�AJ������k��H=)G��'2`�znIF�ې	PL/�4~?	� �ӗ��~Hk8�j���l�c�G� � ǉ��m:cg����r��+�C�}�:�P�6b�3�g� �br˧��=�-�}ݟ�Fy��7� S8�N�r⯝��O�����^djLC�+U����UuK�2Y�9�N>�sXeǚ�/o�_�����jB��~{)��0��m�b�������"J�;����έ�8�Yi�+'����'� A�� �J��ˬ�Y5��T0�3�!~T��F���]��|ۄqrϦ�K}�7��(�Qs\E�"���#�w��,���
@��'����=B���}5撱
�l���ݏh&[Oc�HP�E���hƷ.��v	Mǥtl?����`�J*P%�F�R��qOB��z�#fni-��h�M?��!��hC��X��\��V����E<���`����r�ϔ��#��8���0�}�KhP�j5�7��M�:�Ȫ�X)P���.��S���g%���
�78���2��<�}� y��+��YMU^(����s�s߱�<�������:>z ��)��
Ķǭ��W�A6�wv���Ǧ��^�3��XlxVHYEB    fa00     700���l�~��E����W��X�B��hU�����&�f��*Ix�Uk\���~8�:w�\�3�rZ���&����ƿ;0R�c4.2HJ3r����L���uʷf��#q�M�TI���P��D`�w,�FokZ�����%��TZ���e�{U��sN�PZ���3�RNn|h4��g2�I)z�5"��30���!۠U�M���ϡ��{)!n�:��7���4F�=�o�B����h�3٨�3c���7a$3 �@��֘�Ќ��S�P&b�10-�$o+}�p�D���=���%v
�b����SX��‑�</�D�&w=��Q�lA�G���K�T����t����o�g5lv�>2Mұw�rq����{ɶ��#ǽ4M:2�beLB���hk�T)`��:�t�"�U5o��u]��n)W3����`� ��I��'-��h=}sɫ�����E^��B����s�5Җȫ�^e�Ls=�W؝fބOj^�&��(s<�&�C�.���YDH�/R�N���޵�O�����+W6R����kjrb,'���\wg���z��j�RU2!gEa?ft	���r}�T���rc������R��ܞ�]F�5�Ub����M�����%��N��nż��Sf��,�z+V,ec&t��~b9vS��qR!��Qh3b���T�*��Ŋ~���� k�Ou��OA����Ɏ3��
=�e�tvD���Z8�M?��e�y&��V��+�#ژ��XTB��X;���ո�7��pY��nUc^����A�}����;��2n)�Ѳ���,�Y�J3�Nͻ���v��X"T�X�{�j�I�k��̑|�{
/��$M�]A���^��9�&�f�o\�8�y�e�nu(�y���d(r���ʇ�Ya3�� �Pa��%�Gf�SV
[��E;��Kn�K5�����]�ph�Q%+)X�m�"q�K�k���w�1���ܶ:�ͣ��B�9E�8�i����{E��r �����$�,
���)>�ʃʭ^A��DȡZ�_�i�2H�x��1nP��k5wӏJKx���1�&7����C�7������=�1�`6�A^��ޤW�=�8�[�ޚ`�q"�0��ly$���N��߇u�@9;M�h���Yp�?�ڂW��H&�O��^��꽥�aǃ�7���BÆV����AJ5ji6v�j���k �e�E�A��d�d˪��]�{���V�Ь�uխ�B�4����1C�AH�q:pJPXO�z��#0�EV��'�"1�ϡ�(<��#��]�A3�޺�O�{@V�9-?��Ia����c�*#-�ߌ&�X�lO���w8�X�܃=ܥ�P�ߣᒭ�x�lG	
޻����NO��D��h^u������\��`��l<$'��f����Ȅ�'�g~j���LTuF"3���Gx<����<�\I������x�=FJ��Ȯ����%c�jMY�ղ��C��,�*�X�%B�u�2�[@����ത�2�B�(���>�rf�db1�"�3|3�.Ƙ/kI#\�]�n���:�L�����YӇ�hi:���j�G󜰞������UQ)�O���S�|��o���2�r�#��v�Ou�ʧ�����X��p����2�~Le����F�w�m��M^yg: ���b�������Q� ��#�ф��f�/ƻ���SI� oDv�/�k�	�%��n�<p$�{�
XlxVHYEB    77da     a60D��]s�G�R���yW�z�OR�1O��Q�hdlX�����P� o�e�K����h��B��C���kj�y#A�_�Ny��JN��=�ƯH*��I�2���8 ��{��q�Lg0[naK����<���x�sIFk����D��`�l�Y`���c��E`�oD����ޝOf���韸�J�!�������evɥ��p�+�����,�u��6�tNo�?�_��P�񜉆Cy6
��+����w!�#��-�o	Y�Cz3g[��К�j��oNB΂�]��}|����/��� ��	Z�t^�4/��on_F��������7`�G�ӵ ���yT�ɇ�p^k���(8R#Q�j����!�m/�~5�*UU�1K�|��dx�d.�U�pr�8�s�Z}�S���+�O���z�8�"!����M�u�+�;]J���<�r�,�%3u%�BT��3�)>b�&y��- w@i�y�̖pq��Z��/�-�G�.�S)��Hl�Գ�~�X~���qĈ�`�������}�5�Y�CG�3h� #�Yv�N�5jD�MXl��u7
�Ng�~P�`=d-S�:����_*u�a\���[?����Bó��~s�kcʲ'U�YL̿EG�AR)��<�1���.l[���En�<��`rےd�ะ*d��YIp���5H0v�s'r����XG��1'�^�?����%%K-#�?-���3zJz���/�ǔ�b�� E���n[  )���jn_��}��/�\���p���B�o�؇(��;��_�,������5N;k�T5xCd�k��_�_IM�[�Q_oW4��T��f5k0��A�_gj�7j<�;�X��o��Ik��ʻ<���`��`/,��O�������tL���uQzh9��!���+Kۯb�t�[	�����Vٴ��Ñ��"�RL�L-O�Wp��{F�۟ʤ�B��1�u�� �����>����\��H/��>*��>�x��ȉ�矝�=�g������[L�����^NV�M���6�=y�k���;x����ƭ
�<�"y��G7f�C\�/46s9ϊk:De��<z�0�Ȫ�o,�2<zp�D�Mұ�22�U-"�w�.�Q"J���y��K�]��
��p��N��^��JAN���65s����`q�G�2M $SH	�LO�D���l���u���JGB��t43���ތ�ܤ&��՗�֟�v{�-H�T�T����jL����O�Q�i�K������F'x�@�&�\*
}�p1 ,�� �<>���V���+���RNL�/�KOv��4V�Q���ޢ�c�?�;��	��r��0��$�O�]�"{�r	����y-�eL᫷�{M�fo�U�N#3��$Sw3�O���m(e7�O���f��i�������A0��$(:�r)���!�է�3S�I�y­��(S-L����U�b/�7k�.=�i=#,^���e���.70�3�W���o�t5����������c8�sh���e=��A�W��cf:�a�b�qĵ�:���r"c�v�Ҭ��N�4I�&��k�cr�Z'�h_=0�g;+�A�� �_����;�g�=�9����FX�eFrڝ|�P0S��M8ka0๶
/6/��ɫ�J?+�73��h�S㤄�4���~�O�,M�5j�${"��訐�8��g��}!�m��֝��x�:4�I+&�_�RM�����bjgh<�7�^�z�kh��>th�~f��*�������$x�������ݯ�~)7��V�3�	'�',}��W��Ʃ�d����K��Ǵ�p�I)!;�Z!=k�\ ���)��§��"�IA��\/��
` :��w����KC�\G����<��c�������F��g������W�����&b�d�� �j���P����p˗P���zjq@��.S�}M��n����������W�-���3���unޔ�
�}���I�;ē��
��ZXjE;� I��ѵ���;��E� �kR|���b����:�y�t���z���B�{�6w���%���iXF{�����>ʀ4"�[�0e�����/��q��ns������33m�/}#��]�kv�d=�bfg���GF��0ӯѥ�y��=�b�v�L^E-*哛x���aIl5�}��������v7����i+�Iw��DEȑ�zx�f����Z)�8NL����m:�!�FH�cp7yB�,����N����-uM�-�T�F\`Ȓ��� ��U�1��PuI����*8I(~��Ѵ�I7�ڴ �Y]�h�0׳wiv~�6R]�4?�p�A����6���)�1P���Z���Θ���|p�M���W�f���{^`T��~��ꎟ���Uf�t\��z��S?�H�r!���Z,��)�������VE�'�����}B4�S��s�)a��HT��:�R��.�S�:��`rq��ȵԼ��(6yB���'w�U����&V=��{��n� G��G9WW/��[�j'���˔S�+Ɯ�rI 4�,b=�_���J�	�
o�JMv4.b����坑�fn��pҸ�E��q3� ��$-�FӭC=