XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6�7�)�8wݗ���Q�X���^��N���_>b��+c���r�@4g01B��g b9�Hm�ԟ��Rg?���cv��4�E�)��F�^��g�ɮ�Ծi�j�����)Ђ"'�l�Х��]u�p(����\�3�+۶���q� r���U�]y=a�Ʊ1��8��g3;���ܡ��{�x��)�j���or��筅��d�`�j���?a�M��I.���ꣳ�W�&̘0�4�5��>����g��������~
k����x-�O�5�?�qP�G�_����#fJ���U�\�ZP����jIS�S{�YZ6��u��a:X�P�� �g��k���u�Iӯ+���°�*T6ۊrq�ˆ}�f9{�
�GÌ��9�@���@�'�l)��/�$�39���_��1���F��~���dJ�fD��s�C\�ْ��Ӡ�S
aRF�4����t~�sq�]'��kM+wg|_���*�M�@}����ґ#,�ۚ`N���C��Z�n�����8z��~%�rL��-�Q����X�Q�b�2U�[B(a�������v�$?A��x�񷥆ucE_}&_d��2_��5h��=�(!K%'�ЃP���<P��Q��=��E%��3�WLN�u��Լ�Kޗ~s�M�W�t��?B-1��x��S�e""2�_6���pFou��	I'/��sڤ�u>c"��Rjuݯ����}�+�F�o}f�&D��w�lM��Ⱥ����XlxVHYEB    fa00    2030P�����)Y���K�^,-ɸ	��Z�N�ar;'h�ƜY���Ŕ`;x�r��v'�P��29*v�mW�\[k��s	�r�Tw�9s,�$��5��������!jg�b��*��9u<�3{!^��O \8n7*ɶ�]g���A�eE� ��@^�:��#T�({�ǝ�M��$?
�46�P,�8���/�(��l6��H����V���P��c�^
k����c��D@4�|��+u��V
�2�ɮ�3��"�����V�1	|-W�@n��f�o��]y��f�>����v�MiίdT�B�xhXl��skeem6��я�.{�f��[���,DdH-���2i �B��>�4&���v�nK�x��{���N�W6\�x��c�r}�:,K��n̸�R�o�������F�9�o�����a�1�����8��Y� ���i�Ťe5����6E�WtM'��EF��8���)�<�h?��a�����������@�d��e�
�cRa�j��M��:���.�?	�q*^r1AFa��lW�G	񖠚�IO+Bk��\\<Z�ł<����F�8v�~r�/V�4Kx"TMH��������:�?��ގ|>�J���E\O���*����C����V��k^�*�3ʹ�����[?������!ʻ�{˺H��X��K��&�6iE�I��ߒJ;k:�����2)ؤ�nW�N������k�)c�ɉ�[-� .�Ô)a,��	gզ�;*�
�%R���tS��;�����,���8x(��o&�_�]�M�
69�����ĺ�����˜f3y{�ތ"������o3).+�����*�@�a����w؏^��-K�!�v�ڈ�%at�	W��RaP�~}�}���d�-�d5�}��^T?�A�H���=���xf���f�5���rq�xU���ް�C����6NU/{����a'��S��]�������oq�m	a���Q_"=T���}[N���������OH����K��0��"Ó��b�mR��GTu��/����Qn��G~��ĸ%��3�ĘŌV��0��N��Flu����B�~�Q�ѧL=r�m��j�.@� �ĢBjg���MS���ˠ.�\�]ȡh���e�����
��O��y���xa����w�.�{R�������|��l���ٜ���lO2:,�d
^�;3��cv��}T�옘/���in�	р����Kg������7��>���I#����a<`[���T�S���p%%j3ٮנq���'�����M�wrwp0�'�S�� �Bn���� �����` L>�|��"+Kzs�}=d~v�.4
SNs��i(��~J�'[���j;7����!�>����o�ë����6�^�Զ����/�p����ʠ�"Dl��H��.�J�����P�$�{���Ď�M�Y_m�q���(��Wg
�#� ,�s���d6J�A����c�D�+�7�!#��CHٝl���_��tP�<-�~����k*&���Ы$��\�M�i���L�9�|i��~�Haڍ��ˣ�le���a㌽�R�Xɳr��Q�(������_��x���_�`v���x�wkXb��%Q���N4�K3a�ΐ� '�����mK���9�zm�2%��Y�])��D$�|��WH��#3xZ��C�/�^�.Y� �7�	����L��wf��41d��!�Ll�h�q��U��T�4#���A#1�#��(t�9�jZ6���Զ����kPidb�j|�r��Z�����W��k�p{G���ۇ�Tr����X$�I�i��0�5�~�~��cC���!�l��I}ă����G�h7��W2�V�so9U�@.]Vy������U��0��p���T:zҜ|���O֌ f���;� m�3<|�k� ��w�b�C��u}�]�>��n5X������]�t-�z$b�hyꠄ�:�G��S0�i�7sɳK�>�*��%z>��o���d�0�����+@e����T@����qS��r�[L�%�`=%���6�4�T�V��-�M��h]��JixKS&��G4�*Kju�}���.3;���@��)��d��X�����6LF �okp�3U|�����|�z;��)�%R���L{دx�Y�J��Ǘ����3F�_ʃ�S��$�G���H���3t���f��H���Њ!��M
���:��౾r��+%$G������Әp����X@fq1�>���)
GL�`���5gq�.��!ۥST�b)�g�ڠ:���aW�Iz$�L|��gvI��8l�r��Aj`	��i[>���7�x��cC@�5�s !�f!��=jz�3���3z�Oe�@��$J�xC�6f�)׻hC��URsy��D�FH\8y��o�zU���'s������o�,m;�!��֡)g�����ìl�=��S�����;���D{ �8�º�[vyҸ����X g=ڌ��6�T�VUm��\i]VUG���HӸ�Q�1����Y��m��(�k��- ���,�	�,��� }�(Z
� D�ȼ�E�,xHf~e���9�e�A.�g��%9�ב�HN}j��ӝ���]A��N�s�R���["�{T��m�b�ߞ&@c}p��CK�3�y��\>�=}S.%�T�d���si���k_�NYw�����rQ��BN�i'���X�a�(m����oB����v���n���s�)Dp����[�q(�H��ݴE�\�Q jHQ����P<�BUR��p*���0v.�H 
;�6Up�"
�R3y��'��h�g��<M��uM��Ba.Y��<]�fD�F�q��]+K���F��ߥw�'!�k����EZ�`!�ݸ��F����gH�&�^@>�I��G�6t-ϩ�d���wիMQ�����C�QE���;R���)[�yp�`Y��gn����S1��L>c*ش���=������w�'�:unk�y�Ⓜ�Q�NH�d�ݟ��'|Z�褦�<�fr���w�#���7Lв/���o�C��䩹���� :������\�m�`+t�R �q�ۨLA�ٔ�9�k6�U?e�
Hf�h.���m�	g�Q�Sfx���4����ns�~��7q����ii��%���ݮ�F����������i�=?d�:c���ǖ�p�^��oް@��r�?�r�E^����i��=�fV�״�рm!�"�GY��C�z�g,�LP6W�w�aWv��b�
r�qr)no{��Y�Q����s�*����m�4�X&!�'e�(���Z�Wܳ�)Dq;�*s
���[I��׭�Mu�����Wcc��"�w���MgzTUˑl��H&�n-�v�ެ���Y��Y�}r�:�����1�4P92����2^P4����>6Ϸ�������x2��E�Z�d�*,���^r�c�|O�D�p� �z�k��Q Y��
��9�K��ө��epZ#j׎��M�B���The�Ps�T�YwR.��X����9F$4�Hڧ�T�v��$V4�Ȕ����˗�!h�����������	�>"�>Q�s�V�t�鼤 9J�IR����wY��,�Z%6�
�M��B�����{wl�p؀���w�"�-�_WA�QC�4� ��yf��y��T�Z��Â��V��iMP�u"q����YGњ�)O�H���B탢O�x�����')����艊b�����<�$qVO��%�KV1�aMQ��-�Z��e @(:�g"�)/O���r����&�C>�օ��1����&�0��6T�[�(��]?�*<����p�foE�Z.�mb�v_�a�i��y/�	GؿO��d��\cV�	%�Z��!�V���pG�`g���&>rƧ�8�>&�P�:z�����5�����Z4�awQ�ٳ*(1��N=k��C�i�\��,n����8��lĄ�X�E�m���Z��@�A0^��>.�<z��I{z�r��B��N�ތ6�����Zv�c��x�/ְq4��+W+��O��/ǁ�B�sHnەm�6b��=m�o����T�-�y��|X�_5@�,�ƃ9-�Yt�Q�%�N��4����p�n�N4ゑ&붑��߭{��@�K�; �o�X�E���w� ~O�ރ"�CO�T2�����׫�2T���+�ߤJ�T=bYW8�r�o}��%m����	����y�#*6�'�a�l�9��3�~"z�5�� jp���G�m�Ӝ:���[�K�ť�j��8��"@��ͯ	+��a���X[����0���B���|*^{ݜ�>a��CI˲�Y�8/C���7n�����z[�.��G�E���܁���d^��n#���'�[��@�\��2�lJ�0X/������z�u6��/?�I��s/�*�Xe�����g'���[0uGfal6N5��O҄G�hx��MhDB����Ϳ�to��sf`��&b�$��>NM�����0���Q�y�S��w�6>5{�ih�Ɖ�.���|�-�H�K3���(���Gz�q=3Q�7?l��*{h��k%�F=%N�]Ơ�vZ�*����pg7ɫͅ���s@�ߩ:T�������R1�r9�P�6�Uӈax��u%���A%=�'{�'U�?í
"H�co����ǥ�23�<L�e�u/ArC`�ua�4���.�����)����_i��Q�"~��v�XL��<w;�p�.�h7�$�[����ڙ��l�3Ե6WI/�ne��4�}��s{a>:qڻ��6�;s�?Z ��P�4�e�)Ի�H�q:2�����[���7*Q����-�S)̆�_)�F�-HhCl�/0*&�J������R��l�Z�2y�  k�K1w��E��o꿙UhFϔ:��H��O��� ��>���c�y���	��V�0� �,�m�ບ��u3��ǰ~�p��g3���7N��T�;+�,`5�M\�x}w���;��d/��2dYw��&�(��q�M���pG`]�aR"�݈g�\�>BR���t��Ǎ3`�yy��*�9=�k������'<�kDg���r��ugQz!���{s9H�0���)�*8��X�W�R������"Ǯ�$��%H-A�����9)��P�^��^q�(3�M���%k=�X�B���Y�@x�r�l�����0��z��g �k�t�t4υ�h������`d��%E���>-�,f�m]����a�����JK�pp47��^�;�v<�8莍 �(�
���Wa[(�5\	�I�A�|�D+j�ͪM?�CW9	��R��x*���pүf�-��Ik���&+˱��2�߻�'#Ӓ�z�
.�q�4��JGS���(������sZ������%bi��*�������pib�H�F<b�9�Lע�sݟ�t��j����y�
]����{�=L�Cƍ���@s]w����1N�3Q����7�53�n�a,��=�!�H� R+V`#<Ǳ����3/���� ���"�^�z��o�7��j�O�����q��(�s*�F���R}K�IX�M���ذ�t�E�)X�x/i2�D��J�S�k��/�3�[\�*�Rfd����"����Ϯ_0����n�;D��_K�Φ�+7I�Ll��Ҁ�r�
6v��S���ѧM���j<���ܖ.�vf'�[�|S�qY��� zץ�V�2|���U�T�'�u�z؆՝:c�o��H���b-5��R#�i�H���?LiԹ����g2�6�*0b�D�J� ����L/s��`Zx��A�_j�������]Y2��3�P���u>p��ԯ{(�.gδ���9j$4�x�J7�]rH� b\>��D��ҍ+2�v�C@lѤT6 ;����/���d,��|��klco�QE2m�0�<�b�rmsGZ�r�5�}|e6h�7G�iQsVf����g���νH��I�^�G�ȇ�+(>��Lȭ/�|���D~�p]s��A�742����c8��[BN �����;�QT�5fy�	�n��"��;A��֍��@w��C���󷫽j�a���Hq��9����na�f�Ŷ��@B��
1�h���}*�cA�	s���*2�_yL-��/K��F����x���G�*T�j��ۖ9�H\�M;�w*C[x���ؾ^�zx�6��o��-���W�t-k!lE����0��Pd+���7wC����y��A3PTG�|��dX^���؛4\��󵩐ic�&���5�G�B��OJZ�'���.�1��8�;����!��<�����/�z��? ��2�g�Ծ@�UƁwx��R�0�r �!�Y�l}�q�<��I���Oا&�$be4^�ENnS��$^E��U	͙�E`��>f���ه�y�.Cf2v�>���$���w��=X�<�=S,�mx+�@�������8S0���3��꺷����џ�(菭F�X�*��L���pJ�V ^}y��#�Y@��y�Ɨ�)i��� E��9]B�\lc�g�A���10��"�V���h��G��L4�O-mA {�7�@Zm����|k��'�؟_RM<�	5y%�<�e�kQ�(�à�����,�$�M�hg8{|f��ܫ)Ņ��V0�6�X^I�N_Yq�������Ol{��̾A(�s��Ɔ�tݲ;�ё����b���N`*������[��Z�°[ۮ�7+Q2H�!]l��7��[����@����<$5&9�XV���b�{u�����XM���x%��_�?5�?��8K.U�X���17A$Q��04N~gvzA'����C�;눮
���m����$7��ױ�"-rW����=���/TJL�6I�\|��gvH�Y��Ld���X5p�4�۠�{��
��Ѯ"JG�ީlۚ�R0�����k�MZ�Y5h����,�S�U{��#�F��:*=�o3h���m��
��bʨ�^�ӈ�x ɂ?n�4�f���¾&�w��!Cq�����lkK��![2�����V|;'t�q�Bx9�b�H߲7Z��W�'x=���HQ�xp�*�3�Cw8e$<�f�!I�O[~�9�2~��u��h����|�<�~���p����{@�sx3�E�������������6�u�L�Cػ�a}�Wm��jr������6����UܝRT�9�ݤ��q_њn���p�����?Э���"���O�QTu[�d�h��Ou~���se�?u��=:�R������	l�J���:��%@G�@����=: ���P��Ͷ	�e����%�r�x����ԓ���t�Ĉ���(�����	��b��e�hĀ�x��61@��m�����XB�v��E��3&,hSQ(fD2�v �8ȍ#�L�QI�������j~�.�ܳ��
G�##��
J�ɱe��M�L�S�s��P �9�;��d�決P�V-��=t������l̺~�*	���?{u!5?��b�7�^7es���_t(ۗ�"�L�1f7��b���|I�[�$�o��|(;Ɖ���)�x�I_İ&J��AXJ{ڦ#��[l@�!	��c�H���]�3����ldg�`�� ؆�_�h뽘'"�qhiLz*"�!O���� ɵ�4�oa�p�������m�E�Rw������v�ރ��,�^:�s��W��M������X�S�M)b���O�v6�$-��Y$,�jtmƫ�Qg+�~�㿙F�A*W/�����άR�l6=�?�� (@���Ȍ[t�IA�{eV�M�֧A��q�Z���CV�~�6Ci�,G����NkCQ�V���d��jl*y.��E�N�}n(���l _7��������=C�v���q��w�`�w����aF�-��<�t49�+��E�fxH	��W�U[^�#�;�n�ڗ@��a�K�p��}�8}����+|�C�a@M��#hը�O���N0�{���.���Y����o��y�<ю���75�`�����C�l
��y���㌚~�ֶk"/b�=D�/e�F�&�2��3N.w�ˢp_��xFرw�2�rTzRʡ��u�Y���UI��	ǹn1�,�S"�XlxVHYEB    9620     d70o?��sڧ~`71W�2�Z���T�&�2� �1�)#3������߱V3���3���0��o�+��V�z�e��:F�?]�o,�g��E
՜�Eڿ?3 �E�1`�ߤ�5j`�*�ORe�*�r��4A��&�.:x|yW�.]�f:���K
��U}��"e����IG`���*R�6�jV�<��+��]XNV}i�wpUi6�y*�"�8���ov���j}"����i��5�C#���2]i�^��I��"W�^sģz���sߢg�|��s��Q�	s�m��`�Ȝ�L��C�]��m�J���`�����+8��d�Gq��ZRN�N�lFyZ��4p�Y�u�IэꨳE�j �����K����|�f�@&�	t�}a�gրov q���N��.֩p%�Jq˯�A5���@�W��l#��Fǒ��%mc��
Hҧl�7Zi����Bc�*픺r���R3���9��=h̻y%,�������M���,Q�k�"E�N�x�u�Rfʺ{���ru��^Q��$,@˷����(ȺM��[��Hg���Ж��<.y�B�XƋAi�*"`�#�;�bAЉ@�i��-��[�&�rW]�P����m�α���ؗ�;�(꺇�Aa<��Xb�ɹ�Q�\�
k��<����<�`�o�K�C�Τj����)3g6�>��$���n�W����
}��.c�n�yx�����|Du���#��c�F����&��My.+{�&�ȑΠ�L��w^L���[Xc�U���ޕ���=+�Yd����~8�ѲD��v�ŕl���l���>N5C��<�8ٺ��
�V'�Y��jICB]k}t���Q�3�J������5��b#G~�̆󉧜�����p�u%���"�`>nȟ�	����'"�R�K�3;i?o�F#Y^?f�2�>���1"7���gm��,3��4艷D���.Nk�S��@|��U�{ㅩ�$��>N,bI<�`��ߕ�d��Z�H#_1��ɐ��|0
�V=�� ���Lֵ�|LƅH+b|XLdR,����2h	�8�h�Q��i?ˡlN2@ҩeC�d�zi�DT-<?�J��@+����]W0>{�BʏsAO�MM����E�>�wy���D:]��ٳ0�j�Z]u�1�,Ot[���L߼���Y�)\�t wP/J����n�{B ,�����n² ���Oa�D���Ip� Z�Lf&������K��=@O�h���.`Y�:]��չ|v�%%��@)���,�Z�QqOq�Q�)sv��ª��y�aH���ұ�(��-oM��T�;l �WA��s�pPoo1샋|�,*��K`�_�,?��p"8-���Τޭߋ8,䕱�.y@sI��<���U�<�4I;� ݅���,����� zb'���2c���O<bY��=���%���(�����������<xκt��O��& O ���1 i�� Î��2G�+	YG����0��b~O����-��&��d�@��{Q��')p�x[��3;����%��Le�M_ܚ�`��T�{��������R��h����%� l�=�@UJF����M�Yg�&��(�:��eR8���+��\�<�rYB��0�y�$<��L��P�=�zt�Ϭu�+=ȚHҵf���+yqٺ\��ۑ��=`�k��j΅*���zi�h���Ɇ�y�n�Av}� �����tg�N/��*�4RP/��Bc�\E©�־[</��e�D���/��B��x�e(�7�"��穷T��~R�a�)���s�)�Ƶw�B��<_i�G�C��ߑ'�7gS�!�:X|���y�,b?W�BS\��(�A:�bFBmަR\
�vD�����<�*d[�{��Z��y�i��{�\�j~�>Ö�x�h�Q��TX,�$��"�� ���s�d;�t��ĸ''��. ���K���6��˲�pGD\n�����Yjs��M�8�>�}�5���lmgG�@Jj؞�Q7D5� ��]��w_����\|i�+9e'掴�D�q[���=:~*�8T y�� ���T��<��YU�L8���k�c�2�kn-4�m\T��<~k#��k��I�6�� 䳆�����Yd}h�t���Rb�6V�8����
�w��p�Z��^������x�T!"�r@�X�ύ�mj��^�E���������gױ��v�K�m��_?�K&He>���hm���{��ત��z��Z������^ι<�����Y'��7�L�Ŗ�5F8�R��v��tm�i�\F7RP�?�*U�<��'QG�m��c ��C�[m�<�;����%Z�L���j���&W�p�އy�R)9~č��NO�۲9J_c\5�!��Z�lT��{�"�]�k��$��jfr�8'R��,��(�u��IDBk�E8/C�w��'��N�[�����;��&��ں�p�v̏��#]d������7<��L��i�C^^�?���Ds��:h�}~����D� �w�8� ?&��+�oRE��gj'��"��%sX�―��h������G��<v{���̓/)G3�'��ҠSq�̍��*=��N^ɩ�ׇ?����ɬ��C�v=p�8t��1����3"`
WN��0^�I�zd�R7���U��}��]OȌo�Y��R&����Al2� �#�D#tVbV��hU�ˢX/j��{�4<>�5��X���?�*w�����16��8�u�SJ�L�RM�)���`�N9�6Nn4b����b �/�Ptk��{�@L���R���E<���I����+�M��%c$Ԑ}��A�g�s�)'�xX���F�?���x�4�X�����dHq�j?E�t���) #�'���F\�6R
n���D-��Lc�!L�~h̋R�B4�5l���C1uҬBGb�!�Ok�����"1r�*�ֲ���@?���9)+�S���J�/����$zW�0��
ſ�5���.�᭼���A��a���k�/H�N�4�#P�_iZ�6�u�#I^�U��E�D��a��+#M)����V��Q�3�%d���y	���!xK�f����	B*dO�V��$�Ӓ͝-T[��)6;Xi,]�/�<��a��?T�8���>U63��W��'�1Ix����a���o���9
d_`e�y�J��T�Z�x�Bp<*q|�� ��ې���z�Q��U(�%�"MY���|�#����[+t��W<�\�٧:]�OI�����	�\�qkc��@�c��a���_�%�����"�O��է����y�&�iv7�6E��k`6ʴ��]���ܰ�|T��Ȯ̞-��,IT�L��}e�AU�$����#��^����`��_'�%��T��Y!�(��{��r