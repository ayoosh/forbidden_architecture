XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����A�L�x�]��]�g=B�|O����mt�W�G|�̕K���@�+$��tg��!��#���x��#z�x����(4��F�X (жe@�A2rS���b@8r�ox�X����<]+ Wp��^��1�@O��U��'�QJ�X��yqR���+	o��Ir���b#���ԛ�ݰE%F=sB�y�~��/o~�&O^i���#c�-��s�}��Ȭ�jf��>�b��yo�~������?,���lf����NX��c�g�vB+�8Y4a�z*�C��S�a�c�D�>���OP�^^��P�oAcw>��ܒ�8o�P�d�ZC�9cS��c��ͯx�i@�2��?W������	.�������t�<�S��l�x3��䯭�~�W�zy]��k���oc῁Tf�^^"I/���&�T�GJ'}d11���8O���D�fYI@(���7��ES�'�@X;Ny�F#��+�q�#�(Gq?�V�Xw�T���2��(��N�|�����p�*�W$���`)h�;���'��"��OZxw�G]�e���ÙK�K�d��=*09WV�����3�}7cJ�i���j0؃�u~-��!}��:n}K�&_Aw"�	�u���r[�}9qŹ�Pռ���������sس:�(bk�3�ݬ>{����qM��P��� SG%�`�ԍtA9	�u�Rn�F��4�+����7�]˧'�׏���GS묜;�Tz��5}��?c�P.���e�~q�w�Nm��᧟,��]XlxVHYEB    3042     c80"Ri��U(`�4��î��;�k��������0[�h��S�I3��E@�ex\/��i����A�2\���#o	P�{h���<�a��w�^���+^p<',=�B�']���Y�<��+�-S�w���t(�S?R�?���2n���RgYc���]��\I@(,��&��.�6�$֛�T���/u��Q��g�_���#D��-�g19'�:���� jm�&�1���c�p"!̗�� ���l	;aMs>��5s�3r���b.'ȩizL�L��Lg.�7ה	z�����@@M�zzZJ�B�c� � �|+.LX�����y�.�Z����*�7�Z�A�D���?�v'���(�Ŀ��,��;h`����j��Fh�E�̯����vo���@�~d�o?u6���٭�v�ǥG?��ISI��B��씉�B���2Mg���] u��R�nm�l�`�?t���6���q�#��n�����C�����H��f�I�b}1P��i��Yp�%E��xFX�4!��k�s�����"X&'J�'����f�.��a�J!�� �q͙�Ro�l���w���P�0�7����s�h��hG��rμ�Y׿�Ȉ�W��!tDP���HIw�%%������(�0��p0b%�㒀E]�7�Yc��{�|[�<�ێ�(,1�0���V��,hT��~�ޛ�����z���M�T��3�bNsz�OGӷ7���[��z�m%p��<��u�kn��JD�jeq�C��X�4q#.E;�?��y���o�_����ɕj!�!W��<w#�`9�W��~Oχ~<��GHQMV�9d�x��w�-8ب��<0��b�	A���}':&��s��E�R�=O�i ��$!���6٦�<N;c}
�\�&�K���Gw]2x/�uX98�G3�=�����Qk{ԔL���gwxub�n��J��T���w��d�����
���[S�O�,|��#�
��<UpX�	}����fm}��A���R{9tX���7::<T	��ֽU7��KF�lKL��6�-z~c/��v\;�4��Ȟ�
d&�
mJ`+����=��wZ����=P&����	��#u������g@S��Rd�!������m I�J���j�(�P�`f��})k����`E���������-U����j�$5qK������W�Xj�f	Z���v�4�Ϥo$���G0�`���$VX�}U��=T0f3���֣�dr�q�2,����ƍ����Y� ��b�vNW�	�,�e\�~S��!�-�k���y��K�}����%�xP��_���c`�xm�¡�ZĬ�1�L%� r#�D�T?����k��c�zTo;���L^���������2��N���UTo�) �g���.��y�?Og�3�(�W(���n���;Ӫ�<���B�:��U�I�e%i��9��0^�K<�E�9�I�4�{�Ű�/:)ﻋ^�7pF"QD��i�D�ba�1A�u���Kf��ލ183�����xȧ�b��p>Eͦ������h��-�q*&�m��g�m�g�},��VB���<U�1d���>�r�i{�W�_��
K]�6tq>� O{���(�j�!Li&��J��Of{"�Q�4z���ߌn��m�<i��fh���?�S5(ql2��ےSV�����F�pg��	��фJ�O�Dz��nQ.����P/At�.t���ޟ�̪G���V'{ų��~ͭ�%V����M���1#��Cϙ�w�*�źS}�2gГ�E���{P�H��ȓkB�ߥ���������y�>}�n�[�1q�}
��U�5��l޳R�.t��o�E2k��|�k�UʛU��v��uE��1���$
��ؘ�8�,��l�	���J�sҼ��Ol�	P��w���_K�m��1r�]�a^�^@�������Y�=~�aWDu�_���q�m�E
�bȳ���W_��B��N���th2�}[SH�s�,�h1�yJ����P�KɻN��x�m��?�T����AV8�� a��5ix�xN��>�齜��(f����\�@�'��/�k�̯�ۣ��Hp��Q;
��b�'aQ�uJ�N�7~a���>��g�ռON�:�;c(S�0�h�qĨ_��M!M�g���#I�\ΰ�/fj�-��i�hq��pƕ;�;��S�[�6��V9��Vf*A���-YE�ye���C�t}-��a�)�0�mݨR���E���Q@����֦]�fW��0g�v����mj� �4B���b4 �E
��d*n_`n ���kJ��N���#��gjt��k�}�a��C�k��a�+�����m_Y���9�5����k �����Cg��8)�\q7�ɻ��`�@�h��R���B��b����zUd��fgu.C+v7�'t�?%��e������\Ʌ:10_־htj��G�:nr�n=���.���L�r�|`��'�(j��:]8�iC��(.}����-w�Ł0^��2�PLB� �n�=6��/?���u
��번��+�3��?-��8:0�������K0":9�b ��O�0�<�|�f�2�s2'�#J|;�2U�xC5����0�$�б5�ȝ��@+[nU��8�؎�r��+sJ�쌌�C���e[��(�ɼ=j7ha�����{��*�8˄�(�N��Q�
M��ɝH_��������`,�����Vd��|�Aߛ���'�f�΂�]C��d�y�17�f��ǝ�n���[[�2L���(��(��I�3�s!1�����B��B��'�@�Ú�[h���O��ڴ�	�l`�yAY~��5����*Yl�H�GR�=�_�?
��i*%�f�[��6�b�?���4�3t������pf�M.��sp��W�B4���E�>?���(Ca����G�����D.���z���H�Oݧ�	�
���6d�EL�)o�y'G�Ե*�v.F���z?``�)G���V�W��܂���B+p-Ffs��`_
s`p�,��635�yC<�9z;��US����w��\gk�9��0LY^d�QZ�)�#D���s����r���@P�1-����V-�G���g���>�#']M���.��$��H��97i��d��,���0� �1����|h