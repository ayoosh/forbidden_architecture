XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����U$�rg���N/�M��'ټ�9�ZF�zq�Lz����R���	%�K���ҿ�n'AB7�:9��?7Ku��-`�_s3LfD�Nr�=�&<Ş�3�B^�N��B�.�
�H�
�����.��yHa�'��ƬȰ퀤�`"�4о�:Apx�KŹ����BW����BMX&��G�0��<�T9����������dI�|�3�ݹv��.�o�57�������i=Լ�e��D�6լ�\��8��/CZ��Ewh�K[$�.
��t��H�<��5s�-����u�X�D` ~����qߐ@ߞ0�}.-��_��g���yQLV�@��ށ�M�>�E*I��O��-0����@��1���yU�/HXy���//f/���E�|�����;OO`�e:4+�,΅
�)9��)�fe�I�c���N�8����s�������/1��JT�F�o$�s�����܂BF�d�S�"�l���_�	5k�Y��m��g��7U��'������5Ͻg5_�4c}*��>w�x�;��n����5d���l+���/v;�MBiK����|G~v�a4��Xj"�DT=�}T�f0�D݌����9�����f��|�_�Qd��6tֺ�r����Gk��E�I�Ҡ�`�_2|�[�m�9e���kIuq��|���ʧ���v�:#őr�Y��� l�f���8���')�Uft5�(k1ـV-�t6��`�av���&�Ӈ�ì pı�=|���.Q_�XlxVHYEB    2e55     b00�E�?]���dᵁ-�Ϫ7�9h��Q
�N!3;�墈�l�K�-F�~wp��$801��zw���t���vs�?�˜!�dR���)|��ꈟ�4�=y "k�������M�؆�V�$ԟ�B�~�޶�|��� �����[6�s�/�{k~���`h�=1k.�cwKL��<����.��̭X��pܖ/���7#@�������1�K����(S7�E�c�*\�F�������=��Y�!�ă���?�7�D�Ȃ�+X:��Z.	D�f/K�%YTJ����ƦY��t00){��Wی-��Ix�	��Ut��Ea~�=���Y�	�4������|�:s������KO����=K��'��êR�sea��C�O����=C�g��z��R�v	V8�Qn�$ +��/�-:(��)�X�g(%�ѡQ�N߯=�r�,=70ٓ��Ĉ���%�q4S+�_�vr�\�NZ��>Z��d1$�i�>�.��_"��=��'-�ʩ�Uc%�@G�tw��7��;�]�2�_�]P��u*���F�jT�3Z{5E6���>T��n�`��5�Q^鏯I��0nǬ���a\�G}�:�^�|�� c�Hja�����G`��p��C�,O�b^�RӮD��&.,H�~o��ם�5�����i#�.,^[�>��/hk��DX�V݈�����P}��NIS�9	�)�/��q�� s��,�%ߪv�-�_�3�i��h=@��eT�S�
�*�+/MX��<��BP�᮹L�IKT�8��`𘐣��-6
"�K�[���@��+�����9�<V��F#X���բI�=�Rp��]S����(�-X�e������G9n/]&{:�)�Z�|{owKY�В#M�ftL�է�q5�,-�FP���#`�R)����P��R�c��hZ9��=����������G`�p>wC�K��F�c��lLZŶ	c�����z�^8���c&�FB2�-w]c�xgu�䅡}(���;�ٯ}���A������ �ʷ�&"���e�u.B#0����� �NQo�,qN��i%�6ƀ�9�^6�"���>c�����ޠV1u�x����j�T�6�3�s��&�r�Cy�_h�Iug���2VQ!%�&�+�С߰����-кN���w�]�~~�)j;�ő�I�ז�4=,5ɥ�p�]�����K�ݛȑ~E��di���^YnX�g�CV�^\��R ��֡����H'ylJ�M�NRS�ńC�;�).��su��"�R�d`�	.���y1Q>�Y\bOۋ����U�}�5n���RO�rdU|TY�y<w�Wq�M�5ֲj�@�`��`�+�o��V^�إ�x�kxhZ�a�n(�����.���eSX�Wi�N�B���H]	�q���:a{7�=K5���FЬ���[���֛�cM�!~��ͫx~T����6��c��q�n���uλ^��i"�0�.�򘵺s��~����=���h&�U�\7��M��|i�`#���^yȏ�^�&,��u�`-�Ŭ��4�qc�_�7u��c��	�RrK��*��h`)l:�9՞	��"��>.���q�:��P����Af�]%�����@}�<���`%�l�O�,�aUڱk���閻�SJ�u�����G����b!�K��
@u��Y������'
i.�W�ѽ�Cp�ݏP	,-�s��
�"�*5���Ƌ�Yi�Qu�`8dYD�N-��N�k/��� �%�u8$��N$Q;��K�Ez��ݧ�@�
��p%h��v�>m�6f�LM}��rA��z���������w63�������0�.8���0Ë�`���6�gR���&���{x��|��S�� *����0�R�B@�PË��:�r1���~*B<�U��=k��Ƙ��w���,�����~���p��V
��D�q�\�l0�ÿ�'�]�{c��8|[6b�Ox���i�C :�D��&����MX�Ä�����Y��v�K�x!�R�����=Wx��z_���ʄ�7 -�Q���G����|��.1ޕ>__��V��+�	�8��s`��������琩��|���a>�����;�%(�@��m;jh������j�c��ƚf�ky�xk���G1�5+7���� RB+MI���DM*Ȉ`��*�3о]v�C�9��5���_�h�&Y�&.��(���J�9�D��������Dt����a����#,DB�Z����ID�_�,�Gl���8���Ӵ�G6�j���z�x7��2L�G�j,����D6V�>7 4��*_�����i�!��ŷ�lu�n��~w�Q;@m��F�Q<��t)��C�'�{���y��慖W��\={����_4��S�"�]��5��6ĉ�P����z1�v���v�_�{u ۖ���W��9�\�]����7���Q`�X�Q�9#�NNN;� ���ۍ�*���w���k���x�\C*�]��E�O����s���z��p�;�S�Ì������6`�p����Z�ڠHEL+�DJ,������U)"�����N㫯~W����_3�J�D�􀖋?`��n�4AH�m��<+��F���; �X��=�|R����ti �u�����+�����9�~���
��^Հ�B�Y`l�@�$]��,K�������O0:D>���⟟��R�ز�h8�e�s<�uf"͵�����G����8 qV��`�!O-�;ډ�O�����#H�t����$�>�6n�gx�