XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ѼmU5Ҋ |�#���_��4�5�\1����j�7���0wG��F�XǮ@�y)"�C��3�"����
}�mvjE:�+Խ5=Sj���E�U U\�Xb��}�Цg
7�7��жMAO��q^:4�ߨ����*`��@P�&͡��/*�uC��sS��h�PW���qq���#��B���g2�����@�n2y\�^���x����x�6�%#ֹ���ra�2�#�> �c�[ξ��Z,{Be̺F��V�Eh��(âp���E���Ϳj��?c�1���j��*�s�i���V�������#�f3)��d��%W�wJL8X������ls��-�\	h'������LA,�a�E5U�"hz�QY��H�B�ġIH}�-�����A,��"A����s?�UF{a��Gڊ��9�o����i�9�v��T�d������{�?���!��+ۊn��\b~JX��)��x*�*T|L좾#
I�{S����'�F��ų����EW��Շ۝.�̻�L�����
���c/��R�|�T.�c_����o�mV�|�v���B3e�g�l�n��d����ف�LXm�z�����XQǥdK�J�2a�3U�q̨�b �-��`5����㯱^xf�ty��K'ԉ��L�l=7����r���:e����-�K�ߓ ��|�r��p+hڟ��O_W�т�D���;!�f�k��zI] Y��%*�5延M�=��,��|�o��}�k��|���XlxVHYEB    b631    1a00���;l���\�1��]D!l:���'B�Vs�<��� �~�]&PSw���Y=6m�q�����3Dl����:����gI�o�_cW6[�d\�̰�
��]�^|���ej/|�feiۡzG���@�w������K�o[�ߟrZ���1��Z�v�K<7��tH8����x�g��*;�L�V�����WA:/7����O/��M��̔�������GD) `>�j�DUH����H]�v�ն��_��)�F�{��+�p��.�S�0�y<\:�s!U a�����i�s<8�>^�k>�?@5'�+v1@^��lo��?��d�y~�q�� �)a!9���3n��R̺����%�"�rq|��RN$,���+�rU����� a�椉��5ru/��X.�fšKR���ڌ��M;��&���,H)F^�E�R\A5�ǜ��q�z㵄k-�e��MDq���/f���6"F1�H�<е�d�Jk�B6�|ԔI�D3o�F����i�2 K�]��I-��<�u����\�������X��;?rW%���UU�ZV{���W� ��;�7rE��_VuAxT���`1 [D6	�NV�/�)7$IC}mFQ�U;xc4��Lo�s�ss��G(k���U�Փᩜ�s�x�(_F^8�����K�KW�;�7��~�M��*ű�ص������9D�>r���P� QI��hUJ�̱���a5%�ʢ�+�BPo�T��-��	y��d����Y�v�p�{0�8r.8ݦqw���Ž8og�Z�b�d�¶�e:���;\��V�(�fan�F���&�����7.��l=z���h�5����R����㙐
W�_�-/!�f6���h�K;�ءjׅ�YL�4.Z�
;��}z���@��!�#�˰hku��f� �j�.���c�Qkr��G���)�!Ft��d�y���	�p�5װ'�"�v�</V9s��s6>�����4]��H�S�ÒdU���nH8�R^HJ'܄@W�n�W�3�F�J����)G �$��w�~%�($�~�$;b���fF=V7�U?Hd�-v�x9{�Z�J=� 1�������B�t�⯳P�@��R~�Y�����ː��������@d5i��D�A_{Tթ2ay 0��e/��\�7On��h6��(��k�S��dp�x�;�*��w	�(\��G�-O���{'xweF]P�����"�+1�t��׀I��JN:�=���-mǮ��~q��,1��qg�������Ƕ�Cb����k�@&�v�۳�;-~=T>p�_ 7G���T�/�z��Hg��ڄM�	�k���Q��s�z�g����Я�w,؉¨�?z��
�_]Y '�0���s�
R/ [�V�*S����i�k[yp�H:�Y�_6D�铙�_'w���M�@V��#��v.�D2���)t9[w�Y$d˭�Y�$~N���,K
�X;�1�Fa���!+���
�'O�~��%�䀷�nc�QDW~���{���ꥍ�cN�-��n{�i�n�p��C.���?d>���2�x�(��u��ZQEvTP���)L)������b9Ƌ�5�L��	)��D�q���8E^��C�"��\�6h<K��:H_ݽ��{dp��H�bF�k���[6�Lq�~[
0�?��9���9�02�Y�^#�ץ���ۜ���ixǐ�7
�2Y��P�)v�,kI��?��SH�k�;D6�LYV�L��5�gCO����@�a����~g"���Z9'dZW=���`R�lo���\�G(Dwu�y�d��@p�п!<����T�c�'MG� �ٕx�V&��`���i�mm�Ãf��4�2��;����!��I���bR=��s((���a�=*�k�y�Ń�Wr�u���}�8J�
2�����V7�W_�ʧV`�8�p�.�1�d��h�����Dz�+ɸ5in(���)�L0_�ÄO��x��xyӕ۠h�(�(hE���1=���Q$2K�?�N`̘cbvq}C�3�$��$i��� 㩪�$�o��)�g�-P8.Oθ�!��$��u��IO���w������e��XKlP]uC2iǕ�Y�z���2��y�����o��m�-EA���͑0�@�Jp�;������㘴�jna3�n��K&������}��K���60���$�߯e��Y�:�����L�?Wӡ(���)`�w^T�2q+i'qy����h4W��O���r���tjC�PEݓh�qYdtE`�c|��c׏���5��l҆	`�:	�\��ύ-��{{ou�u#!`jd���"_h�V׆Xb(�cCmE��^E_����iUvV�1��"�P4f�7E�qM��l�ν?���*�۽E�<��B�&�N�o���i�F)�_�T~���S�~&��ϊ=	�e6���c��W��nf��]I��4q�Axٚ�[��e��޺�i��L��_Tl�/(�Ld6Y�j���yr|>Ǒ�_.�]����)p��ة{D��[o�螆�O}Y&��~?��7��|*���)Z՜_�X{�j1-t&��v1��3�i��eqC�*��RcP�W��Y�w�"QDk������R������U�XO�PNX㜦XzD�s��th�A�\�)� G?#R۴��N5�j�.*�z��s'�ߗ�4�[�ʖ� �9P���(��R�]J��c�s���x��.����B��;��O���F��O��8��z�3'��?Ze��ȇ��l�[��g��V�&^7R->��{�+�3��дz��ə�����R���$��Pby�s��؉3)�}N謗.VAE��ܶ�I�F�#�D��H:F<],�D.F�L�, �=z��ݳ�b9���Р��<��'��	X"���w�6�<���]y�*� [��m8��՟�)��#�p�IV���"�kuU��<j ��(��β��cd�㴅yjCp)���,��-��V������V]<�QNZ(\�n��|+A`��@$u��z����Gt��a���5�F�8̧N֖�.;�F������7��j���`]#�wPaVX�K��� �*�F����D�P+c�D�Ҫ�����(��?q�x��I�R���o�g�	B�1��40�L��)5v=�܄}"
�ȍ4�]1?#Kc.�O��¨�V/W`�~ɮ���'F�atǝ�_DĖ[�q���R���<��`��:�'r�t�U�L	X�:3S��K���7�:�xd�n7[ј���A��Rܙ�n��rM�}����" .`�k�7��9�V�6+���d��%/}8$�I��y�7�d�O���[�7��g�Fj�T�4��u��Q't�됧o�XS�}��08�;h���u}T��Pm�bd���*�1O|��2e>	=s?8�)bT�4JI��6b�"��K�l��nC�^b�J`��?U# �a�C��:\������lvD_V�<__xF��f��n�>�Ԗt�!�U����pftx�6�_�w)M��ne7�H����C�SEi���L���]s�9�k�VwIh(�$DZGfa��/��u��U�u��-�^:��V�Z��&P�"ϺѠ��O�vv-���g������<��o�][��H1�9��M���$i�r2:�~��{ހ����J%k������{�>�-����ӱ�G�</[ζ���#��a6��#f��i�ƴI9��w�ݶё+��N��t`���!Q�^tv�imIuNm1EHVu\	��{���F|t>f��=l��CNn�͖�u-�D����1��h7͠�OAUX��sO~-�h�8De�=3���TU��x��,�HY�K1ez�`��ǁ��-�	|'w20ʯ�FX���Ԩ�v���9���^`��(t��8���Sn�w�d_	P�h{�lQ쵀'��#�|o74�dT< [�&h5̌tA0z6���?��=�Nl%�mU0Lw^妊����|��&(��F2d�wI�������R�@�l��ꞙ�Ց Aq�#��dF���~=��]A�u��+�?.3.h�v�5W,��q��߶�"�_��ѐBR�}���	��/�vM�j�O�]%��� �_*��LX04����,s8�{n�׎�Ƚ�����E���hr�^�Fƃ�^��EG�ƟcE��"�p�mH?I̴���.��#Z�l��}�*��2�z�'��J*�	��U���2t���^��ְ��X��wZM6v��{�6���bk�q�W��v�B��t='l��\բ��B�H����e6��9�2�qOmu �6���K� ��:2ꛮ��|���*,��=x��X�>����.��@�����ƚ ����fԯ��k�c���M1���L������ChwY�-�<�C+Ej��-�5*�f�;� 
�KY� n&(4G��=��k����g����Г$P���Q ��l�~z\7wŞƆ�N]�CW��T:o���tK�t�^ެD��1�z�>h+�����Y7Ŗ��]�r�1'L!VŚ���:u�Ui�5'-�|�~<�7|�)�M(s�"���Y��2�f��<I�k^x
�=�i���n��nh,�0-leݵ�;��B���WP)��Y{��D �t ~���S��S�w"�-"o~�����<J�%<$�:כr9�H�XU�s���3��eM^�����w�8����|++��n��vs��0z�� AP�O��?(�5���-�C�k?�R�"��d��ֺ�c0f�1��q�+�NS)���B\<)�ʺV��%r����AA���>�>�Ї�A(��  o�s���X!�.V�1D!7t���'�$*�7�sY���O��8.�n�������T'�&U�j���ķ�r�����ּiF <_]Gq����B���>Q�xbǒ2��ɷ�*��@+����<E�\�N�mk��B���ߨ��)��"������qt���7�}�M�ڼN��+1h>���­�-�m��;�u�@�t�'+�EXF�8���i�VB�Foޑ��}[@��jI.6*�+>��b�%���ǌ,Ѱ;_ۓ�n�̡�H� �����i)�u�G���X敝ʈ��}GB�3����9��ZFUrOOB�!}����Η���P����>%8&q՝Y%*v�T�;����!�嫂����_�v���C����Q����%��D�f��h�H�}w��_�Ệ��[�,nJ57���r5w��uG��$����AGU�(u�oY��z,�:t��炔��4_�0���-�5�x!�v���pg�i��|#x��)B^��ݟ��s�s��� )$ٹ<ِ#V���j����@��q؝�\�m��{FQA�ߏ�]#�.g�	���"8�,fԢ�Hk`'2�`��� �k ����hr�;Y5� �i�ʟ;&���n���5��)�-��:4-& �	w�j��z�F-��X'���V�K����Fm�$���$���S�q!���b��r����)l�B8)v�^�H|�X� t�V�C����Y]�c'��
V��1r���8��F���I�F��� �Q��aӣ��;���K[��#(�[���iYI��WZ���k�隂�����Ȑ���R�:A�O;6�?{���ea�B5 <�VlE�nmѳn$nof���8�<h���;fFO�Ed���;4�L�/����+9n�x��г�g�������LѦ�z�MeR����#��+�QA\��~dkCf@?���o�C�di\�Ԛ7��a��Sr�ֲd�C�)W���O���j�'�'�DPSSq[����8!��j����KetC�нy/���y�f$\���9�]sT�!�)�ɶҲ�D�#��e>;��x�������ZM �LWX[�����r���f�}i*jt�!06 {��z!�w��2��ӓ@�'��֭��@p�ŕ�
L
��'���Fn �wo�o�$�y�9�N�O�{)�NV�Q��y{��^���!�u�VBtﬆ3�z�_+z�p��X�X����	�m��є2}�_��̷P���"�Z�xB�~lX�^Ahު����!���$L��J�1.Kc[c�V?��\����=,nJ�G]� �wՊC�v�<>L>)�IY��<h���>������.�Y��@�&��9㉗��/@W4��_�B����LWE��"&�$P,K�2-�Ϻ+BuqR&��!6>oH�g�Q�>+���r��x%���0����~��ȕ^
ي�,��uk�z��8���?(�'"��3Z!-*>�2�(d3�m��ʫ�(�2�+�^E&t����/���3.r�&�P���0�jb\�*�!���U ���@��N�?�q����&��kU�e���L�mT��,�������!vK�s�]��mG�D�V��"5��uҌ�H_̃��S{<R���j��{{�ryJ=PW���/i�0/����u���sJ�'�:\�]�U�ߩ�xx���{$�`�<� �C�	8zI��1�sX y�(�.��0�Q��*M��H��?���aM��7��<�	��\��C�ۋ��@����D_s��C����ȫ3ą\�=F!=v-�
��1�H��B���