XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T��;�5�Nv|�זPT�����%qb�֯��y}g�_���L�躷�06�v~�س1F� cb0�=�{�$�����w�u�2������uk�~sbA:}>��pf��5ߨoe�e��2�U+ٵ���� ���g��n8e홙��G�p$è�� �nS`�>Ny�X���S��N/�B�~�l	�͙��ɱ̍�.�Ox���j���B9��[�>�)�90�Jٖ�y��Wt:z+�V;��.�Eqv���h�{-z�$+��V�ے~�>G��1��Ȟ�U�w`�؈�<����M�ks���:e�V�vg�z�"��!2����8������j�P\�x���mN��Kݨ���d�4e��B������ۀB�+x2��5��o-<����Ǳ�pF�ަ�G�
2k���Oyt�uq�z�+��"i��rx�,����,G�E�_群�	8��i3��:!����о��L���p�G��`v)���Ck>Z
���*�z��<hŒI�=Ǽ�XJ�G�t*���G	�ł������aVU�1���2��r9~�\2W�JGs�ɩ��,]2z�y�ҏ��^�0�C���ؤ��7���C��s�vb=���G�<h_J��,�~�m?�g~K;+]�S3�ZXL�rK�W(
'�D��~����| k�.j��[7&�L��u�S��C���q�@ ��b��
d����yp\�ەe��ݬ�O��l E�3s�YP� C��_۽�(fh���g��sg�v�*XlxVHYEB    3519     cb0Dw-=J2��#�h��l�T�%]8��I�����y��3���}=E�JV��Ȥ�s�ߖ*�:y��2�^t,�(B�w6/4L�цg�	�L9۴��<��6�ޏK��`rX������~ҵ��>�n!��EKA�o@�.��'�����-@����Yn����z�G�lg��m>�V�!��>������%���0�y��-���\S����y�#ل�����Ap�[̆
��u�kctx�+m~��V �-G���^���X��	�:9�^Kr���4}��=Y���Fp��-ݢ�V����X#�U����9f�4�?b�x��+Zh��])٦!�Wk��_N�j�ְ���&��ۭ��5����-����9����Q��R#{u��/<����+_!����P�7�*�GbM_�hd�˨�c�}K��AHy��9���}����]ٽ$	��������6U�q}Q(�Z�s��A��8� �Q�������B��q�wȶ�\�8��x.�`�2߱a��4,�D�7r������Ȩ��3�n�%-��䊱}݆�tL']8�Vg�{�� |sN%Ů�<� �6��Q�L�9�h��;�}��cJ�'	�V�N,�ZT���O�+�7F� �Υ���:���Y�P�(�,d�ڿ5VXu�=�����������_�3�r73�N/�.��H���3�L�Vt�pdL~U�K��F��]�ޭ��Us��wt�/י�@�|��V���L��awq*J?��dD�W�k�H��s�������������9�S��Sw�>�أV��/�X�!?���u��$�-��Z�E��$��4�9����?N8^.��Z���
�U�]��L�g@׀^��9���	O�$�Ř'\����o��o�͖z�(5�-*��u3ӌ�-Jt�_q$���8>�H�.Y��+;�Sj2��?n#?���c��%����b����ȣ^�Gh��u��s�xQm˦<�9"���M����I��|�D���B�~U=�[���:{�nO� ��C�`�@l\zC��Aof&~y�)�i2�>ݎ���S�BH�s[}bH��jV� �ٴ��ηK�����$
XQMK]����[w�V���Kq?����S{��m���p�����)Qa��ɔm�AӑZc��SE݇%��Ŗ_�7�R�:�#	`�9P־&��sT�xz��q�ӱuĎхz�}��@�az7�E���n������,��\��(<*�j�ʔ���Z�2�����Ck�H�j\Ą���	�:[���j���|���
t��L��T�����jF��\�&1�I=SY�a1�>��{�����[8�7��{ow���4S��:��������}�.4�s�$�ǟ�����'�`������O�xcܠW�ޣ��X�C����uN�D��W���*�W^�1�� ��д�:2�����}�~��qG"�@��KI�ܜ2K��>���]`���8
�x@g�"�4�� E��N�ch�W` �t����"%7�K���bư��Pl�j~�ۏm��d�~n����`�X�����oL��Gʹ.4ھ*�%�������:��eS������\m���n�a�e$�j��Z5PR�]�p&0	����"��%�X�ޯ«Sd1[�z9q��l��TǱ��w-E�S�ոa^!��hha��8��u9���!'���4w���Ù�*E�߃�}"�*ڐ;���8��ß`:4d���Ff���=�)$P�B�r7�R�L�Vg�u��L��Q� ��n�f�<��B��M�'�A�&����h��Wj����j��A7�Њu*�і���P����	���ez�Rh���U��uf=��/���	V+��]ؾR�<�Ŭx�H�]���e�1�u�<�a�:�D�{��6�9�1��	�U(�C^=x��e�cjv�������BL �X�k{',�R�C���vcL�>��H�7Z�Ҹ]~+0[�b
U�y����t���:�Հ=(�T�4}SzN�	�H�:�h�r��ZԠ�z/�U�Yz�m4�B��{�g�s�
[e=Z:�������u�z����nǾz��(�P���_gŷ��BJs��O�풴���'�6	Fa�3�"Do�*td$Z*���EG�����VM�3L��4��|��>��=�9)�}����}�<�%����"Z��ދ}�3l�<�E�0�(�qZ�)V�9���qۥA�p�����].Bi�8y�W:Q���S��1W��o����=���.�*Op��B�q�5�ոf�|`%0"}�宋��uʋ�	rQ99$:j�
<H����
"S'���É���ٳ^�1)s�p5�d���^�گ��b*	z@�w!��x���Kz[JFYIn֕/#�6���1�<�jv���.cr+�[��뙜:M�vYp��d�s��8?�r��kh�F�q�U�b�D�Ǝl��`�4(��k�����r��K��-,9�&
��mY�M����-��#���R9�:U��!�^?c���~%χ�nҊT)��wD������=�� ��	Hfj��� �/�m�H��<?��|~��[@+:�4ݸ��Z"'X���'6�m���t4�䍎��-��PT��_�,�M1(c-(=x����S�I/�5���C�����3�8���#���g��?���q�C?8����~E[#C<�y�qE�G/����cv>��Sd�i@��;�>&5b�\���Q����W̧#�>��͈s�'�EM�?��e�4m����??/K���O���v��i:������Zˣ{���V[q����a�Qo���G��$줕D�4��7+���J6�$Y�zy%
�L�|�]c*���O���xT]%bT^,���P�} 6��z�-R�p�c}c0{�-ӟ͹�EFڴ�*��j� /F���<��g�� �n��&)H���Dr�O���k�'ٶ���A�`k�q����"��ۊ=pe{a2>�Z��-�sF�1�,��Ǝ�W]�Kj?^��a�i/��\�Y�9p�̠��7./v(%Y5C{�s�N�'O���̾b�#1�7[�����DKd\�q�
>I��OEK��ȡ@nB@��!s ��WP���ܺ�?$w: ��dQ�����u��a���^��'~�b��