XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t�������	v<�����7�k�U~?YoMg�K�.&AU�ܘ���l�8�ӒU�¯������S��� Q��|k���AjU������
X+O��k)E�pe<{����,���30on�Z�P.��jp_�${��u���{��w~Ò	����]6y�j@@ɺR��)Yx����^����hvG�ʩN|^��c����!�~PH�w�1Oi
W��֚v�[NGB���"�꯿��cV	(��V���)��ğ\8�v8`0s�riE�����Q�]�	M�S����ч9ɗ�>7?:Ȫkt�?��y�G���ɐ��}��`a���Bie����j`J�A�L|L�$�#�~^�]��Y�tu��r��p�O��`����mc�Z����O� �g;)�ujRj�[d��
@�`Y-.�s� 
��*�&�ʿ5�Za��c3t��ອ�}�<�5��<ܖ�6��@��^�O��|�t��!�8Wl��aI��Gj�ቮ�߁�0�6��p0lX��\��Mؑ
5�Cu�U8{�SW�s3���=�'����]P7(��x��Խ�4�8߶�����z�"aN�F������\ׂL��b�]���0u�֗M|�?GS��/��H��e~�W�)�
`rO?4�����H��y<���&�x����.sI�,$��ll5o���q�eNN�k�Ǻ������i`��T@�|��!nF�	���5Y�>y��+�T��QA�;4���{�(���M_DǓr3�K'���\i�XlxVHYEB    fa00    2480L�1����l.`gO�2��.,���"t;ܒ�(>{%���:��g�.F,M�~,���4�P��@z��a�����E7򖫢��'G���� ��-j*���3��#�g�2��EL�>��������
V���|�y�U@}�	�Ѥ������������e*�?:Yk������5���;�ʟ&t��m[Ns�����u���.R�>���}����ɂ�-���py�}6��&:"��B>�:��a{4Ic�B��h_�8aq�n6�/�bؘ��<��	�K�,�e�\Q9����5��/2A��rX�Y1�<%o���f
���r��c��o�;.a�#�Lg�&�����H'<RŅŏˉg�y�T�R�H�,��W�88� �������Nh9:b��/����� "���\$�t����C:&�Ե²�: �؋�p����|��Ҷh� ��>�	�*ʢ�g�l��E?�:� %�]�k劤��M(�2~V�����g4K�&{YiT��EQf���yDsW����U�S`���܃���6�De7�)��+*��7�>t-�n" �xJٛ���x 	A �U����P�]��k��ŻEiw�)>&k�L���h�������L��H��},w��Fg3zQ ���p�7�E��g6�SV�N�4X�՗o|Y��
LT	��E-qfB襀y+,�K�~G�1���CU���EJ�� a_l!v�Ms���|Hju�\{D�'���&��ٺ���t��|�Wz���B�ņ$�b�z��|��Yl�~�5����4�G�_1Z'��%�����3��@�_�Tp����7*Y-a�Ts��쎍G�wl�싽���0�E�,��k���������l)̬��%X��iV�X\��(�B����Ţx�k`}CO/�����8��+A��/�Z3b��oꠐ(Z��0�'�-��x����S1#}�Ⱦ��ʼ����Ϫm�{�?�.�M���i� @���r`�C�D���y6]�1U?%��C�gy��-�����3
K"�Y����z���xI�k?vw¼��n��õ����>���u��2��ä�����1��A	e1���*�{ad�6p�l*A���:��D��KG�Y&�옔�sP3�E�s�x���*�<C����w�'�m"`i���������Җ�p�&�t�ő^r;�؜��{�P��F�(�� `j�v\3�I���(L4M7���s�ZD��XS��_Mc6z^�KK�%G-�1%���2bZ�)g�w�!fg��tު��4t}��N���k�"-X& <]�DK��*��;��g���P.�/wѧ�U�V��o,�x���N�{�7w_LW�Ć�d-8��f</�o<���"{�=,`��,�|����l@�햕B龄;�;b�^x�t��-��e1�n�E_9ɜ�N}'r�-���b�K�������L�Pu��|jwP�H)��?&m07���$�0��~Y���N/�Pq�F��c�o?ש��>Yj���`ɮ!��T������Jj�݃&�t��O���)P��=���̜���ӫ���Y��=�L�	ׄ���$��w�=E{�^��� \=���7Y9��\"Z�ۺcA��+3���쯛BH[4�K����{V|��lR�h
t�sr(+I��O<�c��5)��Y>s���2��8ިB�����^:jI���"b��B}�Q7;�M�np��T�'E�qG�0������XvNF�|�y���!����t��
�	��(�<G^�|D0�4H
1�ʾ���ױR���e
�:M�P�F�ͳG3%?�E0!�$�S�����9���~�* �@5�[��+�ƖCN�X{~���v}�2&d�z�0rՓ��`�	n�-vI�!���0�,����-�A�趉t�Ħ��V�mTxr��Mܑ�3�7�ȝ�,l)�.�dZA�
/��ZB�}:��
��8A�suOX�%���u�ǤbǊn�3B�`�*v���y:&�י�$��ӎ��N�K1�˥9�;9����FoG��#����>�[���B�z��G�G\����*���y�c� ?��%�Ml%ܝ��\�R� ����g	���e�"���}o3s�_&�G�ݚ�n1㊥[0�'�XK��Z�3�ת�,����u#�³���/֥!Ґ�*��b@5Y�b�Hmǁ��+)����}�7��K���JF�p�M]:U��A�ܬ�&Ff\u!�>�P	=��Fi1��S Ib��HU�%n�B��EO�]���[���m��fќ�f�bRS��|�ߙ�t]����}�F��8g���O�1o�e�����XV�
|�^P������B�W
*���Wػce-��b�A�~Ϯ��ʾ� "@�K����nVʾ� ��`e�CNxd�w�%R7D/�z�k�	�^<��s&��o�:r�V��������"��&+��-e& B<�\����Ԗ��YZ�D�:�:��k��T��yL�]���/1Pg��%�k����CNS��\�JG ��3�:Hٵ&�L��o_ؗs���"kq�Q����DN���'
2�\訿�/����g�q(�c��Esl�>����B�L�Qw��D�j�t�Y�v��I���x�N"�?��ȍ��kB��0�!�.	�\,	��3�<�W`��j���!�Aٗ%���9��8����2"�#)}��T|�Ֆ���v���/����_�V{��M������N5B�9��<�,�r5�%D)pև-Þ"��용y4�_LҸ��:ah��d�N���*UDv`ܣ��
)��DU��x��G�޽��-�o3�`4麿�V]����s�`[\�	������b��G����KX�6��i�[ʲ=�5X�Nmz�O��K�����H�f@u��p�6I)�X_.e+�]��T.`���_��Ik�%*�aBs2���6���gp�Ͽ~JX�AX�wE�2�E\
��  eo�@K��1��.��0��N^	?�{R�
Q�-�i���(�s$_������(ǽ?��`�hD�0tV�����_H1�y
[Q�3k��؉�siO��ԛ�1�׽!]��)��rE�m��a�C� B*l"�e�j�pM�rN�%��Ak"O.[���S���RD����0)����%ê����e6��p��k�g�V��=��ilN&k���T��~u<c��&��y.�YUO��3�&�F�÷�?��(�j�*�Y����V��$'T�\�9����቉�q�a�zm�����6��"� �2ԙ!9�m�HU��vIЄ:1~��t�i����h!�h�M����+�9ʄK�q��*�<����6�ںuM��ٯ�=��c�xVΘ�eY4މ$!X*�+3s$U{�����e��jlТ�_w�tG�f�yp�y5+�"���F�!T��w��� =��>���LDd����U#7��C�s�Fa����_�Ư��!q�ˎ�Q�?n$W��]�_�9�$��Ԥ]uy�V���������u:$��FK�>�x\�{b�2�����H�>-�Y�����έ�D15F�����6?t�X��-�	�2���Q�~�{nJ�y�j\�
:��p������،�Jw���B�:�|�a���vA1EY+���xBtR�	X�n�{eJ���`�&�a _��n�����p4(�Wq��,,�g6��@Z���鵳��tI�\��G�{-$F�¹��h���L`@n�^�mm���"��W0�_�J��x\�1zp3e�ĭ��ڮ\����r8�=H��;��t�d�r�.�.9N���S�y)��F!�dMU����W���o��Ĭ\����
b�U��DXءKq7��.�J��ˢc�9g��M�r�B/_^�B���W���w�2̖m@�'!�r�=Ÿb�I@?N�fg.�����MNzzB����̉n�3��D+B昖�=^x3e��	��j�iNP@�8�ǩ#��G�������b����U���YX���� -UY�����Y�F׻D�a�ov����ԗ�M��P�d��yˊr�6 �������4��N��t�z��eábQ�QF$+�s=������kv��mP|4N��4�F-��C�T�dr����(�����C�O��#�sΚ�TF*đ�2��p�;����$��H`{���C`�jފU�yj�K�熥H�׌���c�	���?+&U�Ŵ�f�`�2B���⁅�	OG�BVV(ґ�Q�,G*G�7��yu��"��V����
��×�P���盳��[p���~ى���W�j��������`���]���^�3����tkI�|QU���9X#}�����|!�zN�S�ʘ9�`O����K��!	��L�H�}�P���)�|s7E��'�h�w�=O��P3n�
�D�e6M�!����<C;|��o��K�~��#1�W�/w�R����9�6KÓ���-&*��
�`��-��i�E�r$��vD��f�*[�@��?���۪��<����?2lrl�B�ǀ�Q�#�l���
�����_#���{�"�HCf[�D���L��#�h�OR�������͜n��^���Df���8j{VK�J����MH�g��.��6l� ���9	8-Q2��u�-��bB��p�M]��>E"� �#J�1�u�]a��+X�\/v�۲�
�t�tSߣyu��y.]�7� 9a(6 Ǩ���$��˄��1���L�@�ʦ֎��Ѡ&�Z��.��8a�7���`.n�Հ������@�q�N:���\A��r�&��A/0�on��nS�*��{���7�|ỷR�d6v�fɿH��w���s�yb�XP&���v\1g� �v�8��%���[����?��,ϣJ��D��lFF5�L��A��_��n��*-od��$�@0�hݒ��P����=.Ь�Q{ӓ��,#{�wh�o�olմG��8{n̒(.䥼ք��37��_����/�*e��Q ��P�?j�1JUx��j�ā �+��ۏ�~2dF#�]�n���<�8���&�׷Հ��~
1��$�GV#�P�G����A���i@<D�VO�)�!&ճ�ZJ��Fb$V?]T��d�P3joCqB#��O��&0횕�K��U�*���`��4�7ȟ��y�0�Z�g.5_�%�x˒��nܼ�1�^S_ϊ����z+s6�١�ZVJ��N�7�=W<Ԝ�̒N�if�S����ܠV_~����r7����P`�>t���sqvi�jsD�*�^8���&���aH�Ka.�����X��4��EY��*�9��1S�\2���D�:$h����!�wV�◛�K��٤����k�*��5�Iup^�
�\����]����8���`#�B9��J��!�&�q0�:lzv��h��M����(P 6Z��Q6������0*�I�x�@�����(o��M�����a^0��L�	�浟f����W�Z�]Y}G��SU���h1+�~f-�a3^KK�"���
.B�t*ּ3�[�v��;	�M���U�ٶ�_����\ۥY�1�����"}��L�ϡ�i0�<&��,؟Ծs�,pTމt�}7��_U�{�ug���}ٗ(Us��w�$s�P���)ü�1jJI�k�BOK3ϳ=�߶��*z�*��,g[���m`�`h)�m�������{���;}--��L=��rNo:�q`�=�e(h�g�zh�7�ppA glH������<V�zձ��WW��+����<����A��a����ܯ|Bv͖���&p(��"0te�piռ��Za�|.���1�ٗÌ�뫔���إY�T���6�R@������0�w�ObKʭ9�����@�Q7����ܥ�(Eʄ�]]օu���b}S�LO 1Z����q��JCY?ۅ#Q�+jXM����\�Ȃ��w̍�z~G2)z�����B�:2���
�q+�Oi���r ي	Џn�PJU�8y��q�&�P�+������Z��T0�8�<չ0��� Q�hQ�}oP"�C�#����4���u���Pjf�q�N��N�����~�:�����XS�;�"��C�	��:-׬��P�M�RfH�h�|_D��kזr��]��P����xnq��e�>[5OB��[8Z��6��6+&�7Pma,���8��#M@V��5�*�%�=t즩��}�{]����xvc�?X����ߎ*�
d�}pt�x~dm�	���sm +�JI�,�{����0]vS�+;��ʒ��9�&B=[��h��ӌ,���B``�%���.���*S-������ض�9[f͵r����i�
Ȇc0�Q���eX2W����ho$���&���ʉ*�(٧�e��.��л 0�	�ȱ��Y��Y_�;P�qѤ���h)C�]lխ�h�����x0�W�Pt�9�'I�Vn+e��O��e���7fɖ���N�l��B
o��. �! �W�Nc�@� ƌ7��)���%�>x[	O WG4i�����o�S74�=�*<��b�W��"٠�J��le���`���"$�ۭ���j��<F��d�Y�D�}�fI�٤��}ٗ��D�7�&�l��%>Ȥ���(�I�
$��CS<�~��	�����aoC����vf�6�T=��l�Ϋ���Z�FF8��N���L��IZ��z��D�8�� �k�p�.6�fn(]��q�#t��DX�]���1{U�4a��pFC���mo�㖚�U��vR�)���D�I��EW��C_�9�=����N�iY���%Zʰ���	gZ��>Jk���ZK󤄡z(2G{�����_���s���@TV(`iv7K�
�����aq��;|B!�^�l��Tj.�=�p;���*��M�[���O�4)��3?�ԟa-itS�е;�f�,)Ӛ��,,o��+�S�Bz�X[���Ѿ�mƺ��i4�9�r�w�Zո��ư���O��D@�E�L�����	�u�\;&�wI��{�4[�s�p0�~(���+��p:F&N,N?z��#�3K@���?L��H��@�#	�j_����4nX�΋�꿀4��&M����G�MW��'g�V+TR��ST2pwwe*�ۀv��r��C{���1iD	̠⠖X�+_7�������s�Db�ȭ`P�>$=G��c�!��dG����QUT�-�bf1mZ8L_1O�t�^X��H�]�=�Gg;�ٛ��d4h��{%�⏺��;��2B���s���f���EŇ����Wo�V���GV)V�������T#ڊ���� �����ލ��:��Gk-nH��w\�Q���6`Muj�>x�,z�z�ϻ�I�Z�e)��n8r^-�G]'xZ5�c���oK�;yrϢ)��n$�X�d5Q�oiJx�6�ZZ;�ߞ����Fe�����y��sқ��>�Թ��=�����%��>c�����~*����fA�KƓ$: �V���L�͝�\0�lVp�����8̿D=>I�a��]��[L�DӜx��A�ɗ��e��,�O����55B�@� �%�,���7th�j���r���=��謫�u�"�J����<�p^s9��t�m8K>�osfK��dt�
5�<�z�X�[��Ėx��a�O�����f�
a�H��ࡲ�R������r�[�QhSf?�i����i�<ƽҩ�k����"�Op�e��Br8k�a�7�9	����v��v;��Wɂ��t{ƕ*�'ŽfV��I[�����JY�Km��AQ�4���	�iz$�� �#0ԢGl�o�����ģ3�������#��^WƋ�)R}겑��Kwwl-"&�,_"<����إ�����g����:WDa��`�#��c�X/���:?{k���v�RZc�)4�m��m=��N��|lq�����B|+=����MG���e�4~]3�oQ�^��L��y�5���do��ϩi
l�W�y�[ѓ�h�R1NJ�}��U��^���Q��Y�=GҍOR��1��T{�_�݇�r,�x��o�%�nW�lC���6U	�n=�:��q�ϡ���/?���$H�x$�S���$$��~�}��t��Z�o0:��ɚgo&� G� ��� �Y�OZ~���hX��S��mi����}��j�`ҁ��b���/V��53��r��]I��K�|�0����OoD��ƣ8J���*y߰�rO�������V�Y;̌C2̅ F#���kxj��)n� ��'��σL������)R��y?\��K�^

,��k"�V�̖�Kqù�H��ʚIB^؄��NSN�#��_#(��AJ6F o�"o1��u&��7�g׉��6�0D��g�$�afy>E�|��k>����Ki�l��-_�혽9{P��G�e$nȗ�pe���KČ+���y�55c˂�V��t�.��G��_SjCS�T��v}Ʒ��-3�߁��$�Ϛ��]�+Pe�7���=A��	���Y|���8ow��y̴�2�)I�|`>Cxl���2J9De�Z6s�>�%����۝�7��&���5��	@��ƀ���]�+��<���<6���q����a�:�3K!~�;��y@-)����A���u�� )�"��<[l��=��/��,�<Am�M�
t'i��bt�C� h���j�:�����jq�����Zpj3�B��R�2�e(��R�Ӳ���4�nC�ɳ��=f�*� �C��Ҕ�M�B˲;b��-_-1d��ɿ5��|F�۾��%�d8F�ϊ�]oP��r.�S�E&���=x��!���aN������b���pc�u�;�!�����@P��߂N���ݦ:�d����|v|�g"PV��o �|wԡO�bz��uQ��,7dX���������^%heT��ua�D1�A�!�����\[���,�j<m�2�>7�ݸ��Hm�ZP����ck*�ա?���'  �L���G,�ɫə]�b�Tv�Oz�0���}�q�������dG�q&�@E��)ʹ]y(�D�AjfƝD������`��<7��X�� ���?���f�a=�F��|��YpB���rOS��� �����F�O�� ����P�$s���=K"*���_E��*�Ai��}���vIC�|��Ǯ����:�8�d&ȃ_��1g��x��N,��XlxVHYEB    9663    1160���ͨ���4��И=޽ io�2�sb'�3|tf��F<�u��fu�G߄X�>h����h�(��-�_�5�^w`-z54c�n�z�o��1Pj\�っ�gX�q���xX��dZ��/�O�A�Ļ��P���&�RB�+7�_m4�<���"���6<�9E��7��$�#	�KR2�����w�u����d�.��	se�H�
����Vh�,���2OT��/���Ҩ�Q����"��q5¸U�$D��d��3]K��GS+۟=�U�X��^ic��{d�� B��lݑ�H�M����,�61t<��R�{/�7�N'�=&ߔ�\�9@�
x6V�����}�vYM��جdF)�e���h�c�T��E_C���:��� "�x�8e��e�� B��Jw0��8 �|�C�6��+���έ�M�4`�L�������I5�������zba��*փ{+/ޘ!�UFeft�z���T���P�{҃U���5�#7M�����/�[{8u� ��5Ný�_�9mƞ�~�V��W68�ӿ��d��D�7��֞�/�r��hw��T8y}�$P!�4п+�*͊
yTI3��^�f�P9t/�E��J?w�����Z��ğ���4-c�O(ת"�5��_N�ǁr}�*m�d����b�����cu���}H�j�	�mW;%X���>�Jۀ�e���#=�D���S'��������8U�i��|I�Z1{ʦD��������yy��ڋk߷�T&�t�R���x�H��LF�?�	Ä� W�i�-}��ت3las�{��9�"����k�-�Zf�����"�k�EQ�M�ͽ���	�\=��Yox�j�C�Y赻<tA@�-�0�w���,[2
D�y�5ˆ��\�P�t=�B�nGs|V�KF���W�1�Ibx[����z�N�0˵�8���DI�N�� ^]ё�K��&��
�����C�Q��qn��T��H1�����X=��[r'���[Yӎ��\�X[� ��������7)z�
� �M�?B�C� {%��O��L�t% ����Et��S5���y��ʚ}o�?vv����ܕ$R���j�+O��!A\t0�b-���κ ����d}����X��"P�CA@�n�m����.�p��6�������v���p@io��)#qĘ�Wd�X����.a$��T�V&9��@C_5G:i2�ʛo����Dp���I�7�\��J1F����Cס��#r�b����^\�XqxQ�(�n�0��F��lF�ź����K���7p)��#���,W���j&]J�6#W��ֻd�E�q�F(����I}5X��&q�|���?��V!�w3�bNH@͵���{�-{�'���u���,� 䪒�:�#d���W8i�+y����\�r�%���kQ�֜���\0���vb��	F*P<f�� V#>b��u_=-�żR���Go�Iwr�_U+bۥ���?̄�/��������cXL�*9��F��m�NZ�7��I����@u�z���5$�4�y���8�{�؞�+y��h[k�a%)�C���U'	x��%<A
��O T�2�w}��?�4Y�Y:��s�{��+,���䬈���
�<�DM�#�bw5�Eog�Hj9�>�׍lgd��|��5��hj�Lkd!-o^	d#Y�>��E���;���l$G������o�=K���W�O�%�_C����g�=�����|�^�?�0�G-���o)#ߐb.��m+�7�2�Z�N�Ih�`)���%���< �S�ʶ�:#�{��7|�	� � �c��/�t��H����5)Ȑ.G����pU#���$J��r�i,Z���w`��Ǧ�&��2��8��պ��F����I�����s�T�AHd<�����I��vlc��[�J� ��c��}�J�L?U�&�OR.�R �'��������~�`Q=����Ͷ�v;,�-�z&/gmLE�[��8��0B��(�y�)}�:B�׸@ĕ�:#T�&�����2��ߵ��F.J�a�4kx���+V�OiqFg�"�yh%�ϫ�zd�H���#��kӷe޸-�ˮ���Ռ���K��noI蘤��O�+��q�U��`��j��l�E��5:M�" ��ΎG(z�(�!��a�����ځL#�p�2!$Z{6�͆f���
�����t恏s^*^Ҭ�y�^w}ԯV/�dh&!T�4Ε.�|�
���%�M��od #l���)w����:�l$xm7�XpB)��ׁ�d"����{w�����)��T�Z[Yw"�l�����g�Zl[����1Ë��ST?!��B�{�/
��p��5����i�@E�
�U>���V̟��$x!*��u��iU��Zg�p���u&^�Na��=���d����P|��[+C�+��>5tq�����+�ǳ\O�7^�F:���5m!Yu�>��%�b��pb���b{�m�	.~{��]�mTl"�5�������V�;o�D�rP�\A�8�A�@	��U���`Z��]]�RdG1�`'�ל��;APG���r���6s�����2�0x�j�H�,�J7�Ըs"]U$�U�dB�c���1a0�uWP!���غ��F}D���QI5=�K`���rorD�6�h�9�u�&��ˌ��w��Q����C�Vi��3	�8��oT�6�FX��x��х�)C��5'
��о7�U��x�4y��(�`*�>ˇG�w+����7y�0d�w<nH��r&dj���8NF������8<�h$�.��� FX�"�ݘռ�����s"E唓�a����y��%��V�����-r��P�m��@����%��<�B�nt��}~�6��8ا�j�����:�s�����c�t�3�8���a��I�KV�Q� ��1�p$ @��A�k<�]�߁��F�=�7pK�O�h��PRV�Wxf�����&Ȗ�;8�/u�چ�W�&���d�n����H��~R=p�h)��%�{,����gBELm�$!A�,'X�{l6��8U#��C�#��ۉ?������t�_��\����شQ��mO�*\�i|m\q�=���6�A:�/J�|k"��^�_���� P��*@Zݿ8O{$=kO��&}�,�Zdo�� L97�E�˯m�������W��N֦��ZW��l���ڷ�춫���'��hϊ�Ձ)F�]@<�'����ۯ�\�~MG��G�|���1"v�c�"{W���/ab����!����3V�Um{����[Vv����� �4�P6~�@�T��͜Ż�^����y�|���չt8hL���<`�Fa�����٦��ۢ.�#F�HX�&^�k�����$�#HұY�����"�t���A�P305�P��g���ޠ�Q�
��Dq�ۃm_���OUq$�jǀ9��9�"8Z���E��K���6�P�>t�Z��Y�]N��~����H:&5�z�gv-��c�ܜ�i������U;k.�J\�8ca|�k+��v^���g7)GV%�)��;���ݷ
�M~������k��-�jf���z<�%��'DK�SK`��r)�/j6�W���(p
���L�ޚ�B�ڹDT�U�L��L"Q8���Nb�Vː�6��_ߋ&�^h��*�7���+0#� �q�^���>-���92vJv��o�٥h>�(��/P7\�lu��º�9 ~f�@�����!9w�����t֕����ql���n\����tƯU���tJz�̆B�k��^}7��x����FzFX��!�1�{ۺ����L�2�;���Ӻ{ �c���#�,>�0�Y{���b���y1��\3���Aw����]�z����1݃XfA+��b�ns�e����2��4��(�ǈ]�6���:�vrO^�ڒ�Gb��{t�>�����; �~�pW�_���:��X�.\1�g��o!"���{Fϼ�9�h �ý�$�k�<� 9X#��޶���	�? OivWI�UA���ݑ�;DЗ�q�i0Ww��-e� �l��B�c�'���@<��������O�c���,�w�fp����PR��dL�xgp�0%![��神�OR\Y9E�������^çU�tʡ.?��׉� �F�O�0�{+�
X���!�j0�]*�ݓh����	9�0���f6.���`zQ��t�''v�����6��L�Td�ߥq)-i1�6V�ƥ�������L��XwżyA�ia�tj�"��N�dU���Ӈ�
ML����I�M�ԁ����(�79�'�x�d&{6 ��2N�z��>a�R��P�0��œ~��_��eHN�Df#u�����A8�d�2�fO