XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|tэ-	��Ұ���5X7���^i ��۫���pV%��E����^P�Ҩ��xȗ�]7��Cr�0�8�6�������r�QE��$X�\:U�=��/�s�
SCxh��L)�TB��`�Ⓠ�Rodh��h�U�h�f ߚl�PH9C�*^��!��x�2�K�A7�׾)�dD]�	w���|�������x�fߋl��(��3d���#��/�T[�$d�T�!����� ���$xJ�J�}���]9�5��d�":��s<ՑM:�*z�9P����)�u���CU�I��3��eJ�uJ���Gvh���ˏ��o� �"�bZ�l�l��$�|�j)<-����݃޷P�VEb��{�N�dC���Ȏ����S�
��c�v�-�{r�a']z�D��2]熳J��nH��?�7|�xp�'J���f����DBw���n�`x(ʣ$zxk�b�E����̪�L��̘�cI%Ov�Q��*�{���i5����"E��c߱|���qh�7V�q�ˀ@��~3m���^���$��=ΐ��_* G���
z� \_���(K�;Mw	����#;�k��l���Dש�D|J�0��Zk1��*��\^�G�S�'���ۚ:
P
�B0���T
��{�½J�騱��mQ�����_5�\5�k�M�mVb��E��g%q �H�"ʿx���Z2*�-9�q4/YS�<����!6 ��*�ݗ�~����	8)d�U{^Fm"�M�<qXlxVHYEB    9747    14e0jh֓5X*�����`��%ax�<}� 5G�v��Mcx���N�Yk&X��=��]$�T9o�F�O���|d�I?p �������{���v�q�O��}E�������B���/[�jL�a�	 .�"r�`״���Ͻ�@sc���Ǳ᠋^l?`R����[�';p������):�&�\��J��F"Az�t�=��]fC��.FI�|h�ܔ���̿d��/�#&��r@fm�?�+b���=�j��>��n�`� �b۱��PZ�"�~X0�9�H�NۮY��}~���Z�װ�k�R_�@DM�)m���R�ev�(��{*n��x�"|Q�J�S! �䳬��\}��Gl��o�@��	�Y y��6�`[Vb���!1C�Q["2���]�V�_BI��6�*� ���lΏ6�+�H-x�6[*���ﭱM�I�/�o�x��n��1ʲ�G�Z�Z���Qw��m{.Eg�ز�t����ưG;[��6��`Z��g��T;.�Tr�����i:gk�
�+]���̦�Y9��Pae���}k�B�,'BH�M	���&k�#�5���1����y�1!G�*�������O^�W�0��ktP��W���|F�F����ȣ�Y�+��i����)&�{\�<\!$�C�����6� 1�ZNN��������ukW)ϊG�Rqo�������r������5�2`���1���F-|�ֻ +A�N�	�~LtO��W����� ����:LE]R��]�&I������׵�@;{��h��!�uz�%$Q��P:�)��v�X;���zf�fO(�hc�q��9Q��m��py�����SIz��	���_��(OGT���]Jـ&����,��:��"c��X4�#�����/}��~�!�V��vohG������w���i$���ͩ|o�DE�慓5�o���Þ.��'[�3c�9�O�Ԛ��&0��~���;2bÎ�s�dJ�]
�'�ۭ��0l�p�+el��{�!$ة��S��V@��Y����k�����p�����{@�>�Ktڗ��M�se��Pl���� 	淃��������8��w���ʣ�S/!"rID�
sW݆�%4~��ѢPU���`���c��:#<�>�ZX�]������}I�%׈u�<8��T�;���6�E��:hL���_���-x�
/=�/��2��x����kp+�}V�;D���i:+k)�tm���(���q���?�S�Me��V$�/����GC��F�]sN�r��r%`��%G%vḢbɫ3�01&�������Z��+�#����8肶9�����3-8��I���g�̯q��T�ey��h�\�G�c�S�r�Xl����(U�+N�Pk��S���m��`l!Җ.k�[ۧ:m:�Wa�(L%e���W��f�vQ�V���仝�����"O�<�܆�4�fa1z�����*-nmE��[J�j���U�V�L��ʯ��|[���Ry|3!��4�n�Di�,,� {$��c�c�8�[��K��h�G�|d�u%92�<-w��]�J*���s��>۠reP'043[�����?��*=�m�W�:�A!�B�u��2IB1
cV��?�B��`����H�NjP��eF��{���<j}�����+��,��b>��Ҿ�v�A���\��ŝ���k�2x� G�QMGh9k+��-B���,�5$Ҏ�,䵚ӷ�S]�屢��B(w�$�'p�9�YB8v�BLOE$��Q�Vf�~����3;V���w�Ϲ!��`� H���ھ?a�`yjl�s��Q͘K�A���a��S���	�1IG��>���q4�⊰;DB�ӷ́�=���ֹ�h�^����񧆞�����~���F��2>�if)Ø�e��Z1A���r�FXJ���1�/wR���P��� -^�����hu���w
��ce�4�$L[ׅ�%��A�3H3Zl�or�~�PK�% wQ��ܧ��a>��,.@�'���]^�T����*���h�s�{�+� {�[��G�S�Z�>%9�&�T0��ߺ����g�$�:��� [��S2C��W�9�y��J_�ē����|�3��2�h��n왕↹8|y���NW����Q�Z�z�&��t�p�;���ĳCP8�Sv|3�
���&�M���WRg�R̭��� �>T�p7V@鼲Z����b���ec���R/eVK�� ��h`���)u��;8���2�y�0T�O[����v����X/��o�)!����	�Ƙ�|Ef�1����=+qd0d�4۽�ֆ��w�wr����bī9t{$�x����j?*9�������H�0Jx�%�j!�V�H9��1�,�����
�Ti�Q�D4A0��>i���rǄ�SLX�=�f���y��5��2�?���W�$Q���\�6:�Q/���R����O�Ih� i�y3��C�m�klc%+~T6k�C:��I�����v��Cc�$�1��~Z��>��P�Sa��C�,U"rΐ"�������O�GR��K�d��r�Ʉ(*�B��4�4'�������x]r����м�_�%o+�E��}s�8����d����oʑ�wo�ϒ�鱷�T��4y H�
�(	ҜPX�W�>��#���\ɠ�g�|�I�eRn�
J��'?�go�����Ƞ[�L{�[�rḪn�.Ā�6��=}�������u�S}d>Q����w]�3�QF��M�����S,�ML�D��_9�3#��H ��	�U��b��)&��Mu�䎂{E�|v�8�?E���yLP"r!�BZ�s��t�����Of<�Ip)��a���`	%�b��l�L���P]�=+J�ZBu��b0F��'k��/�J3�w;��*��>�������L����>ԡ�}G��#�9��>���N��I)+���O�L����kb�wnaG�ξNj߰�.\�oP<�kz��M�����o�eR~��sx�����lQՂB�P�qD)�?3��҂�����"_�4�	�b)�Eq��T�p�瓖��%;�2�H�	��ծwp�"(@��� m��B����Ň�T��q�[h�q� ��K��:�Z�:��]�-,OG�R�	I�r�k|�b�'t_\����a�G��b㤲�{��k�	�:�+!�:Y��d��O�����1�M���:߃SU� $b�ьm@��~�G��fJ8�T}�:V����l�z����ͽ���=>8���K�� j��cO&�����r�j܂��{q����~�'����^n�N�&p���q�� h���$�[eƮ2�Ƣ�Ǒx�i=��@�qШ[��'�?{���a݇d�BA:��G)>�\8/��[����Kj�Z29x]�4 ���$V&'���ܾK6�:��EZ�y"�5�ހ��,,� ��a~�]"f�诠�X`���}?��8S�.%3��^a澢n�o��e'�1.&���rj��S������T˒��n������W�(���L����^6�Pdm�#C�雨4��@�r ��N�giؿ�� ���%�Bk����^-n�.
~�-�
7tk^��c�D'麸����Ī������G�ZT�<��A�?1f�L�s��	�<%�r��<��9\�5�xT�Ԣ�+h��p���%��3���Q���0=�G��k���y�3U��C�5�0$qOG�?�|�poR�{Ʌ�~韵��K�ā(��)�ms�k5�� ��m���*L6w7��p7eOZS�a�[ʤmff!>��K��"��t���w�s��E���c'����J���o{J�jy��
R�"�fd3)\d�ra�֗�IC�~�b;�z�H�9n�ݽ2J�IP_F۴4��C�&8��.2��+2��r�%e=��� ���غ�I���.s��#���3��3��#��`;���q �
���N���=k1o��DX�2,mGI�F�%ˠ9o:��&�*�i�30
,[1 C+\�k)}��o�J]`�Idu\Ge�~~}H�����	)���w��֢����+���r�/��q���Lb�pk��.�/�DwE�l�E����2������/88�.���+�Q�B��/���2ͪY���t��/�
��\=��C߄�󮗘*���;7�{Hcr���C�`N8L;Sⷀ�]8	*��AT̼�v�Q����eZ�ARK``�f�0��K����5�2����Q@�/�*Ca�8aq���T�Q�t:Dٙ�<�7���=h�^�)�ҝ��Kf9�Y<�q��:��b�$�4�����զ�1gv��q!qqwu���n�d�a�F43�(߸id�Ӵ��j��9��m�XŴ7�q�t�i-��rjղ�\�!(h�^��O�����}�m�{� }���;���Ј�>�a�/�bi�+#��I����p��������G$�Ζ=�w��h�7�3��=����:C��ɏ�!iFYY��j�! {��8����vP#�D{x��`���F���Ԍ��C+�;���ݜ�h�ɓ��.MM�ژ�S*�<��x�\ŷj���R�g ��i�����c5�TE0n�ԫ�Ƌ�ΐ��O ��H�kŶ
�����U��6��G���!��rc��mm���\�G#Z�������3|�����J���ݤ�v,�R ��S���nZ���i�4M�P�X	[Y{�$�Q0(��Տ/O�G�s��c{����-���c�+��X����
��S�P���^2�-t	l����˔^��<]+{H���/z!iT$D^����x�R=�Ш���Z&Ε��kEQ������=�vό<�x0H�0UAd9�o�vEr�.��,>��U&p�wH1����F��h�<W�s�лaR߻}�E$f>��;0M�Me�����H+��p
1�j�⪳�3ϰ�����������"�q�S�k���1_�D�y��鳮;U2sH�0�#O�/JY"��qv�+a�6,<HΧ�1�d|u�����dЪ�L���ĥ�����l� fW	��/��Z�Ɗ6�>�/}�Qq'J�v��)����P��H��F�5�����F�]��<�>���.(� ��1��"�}٫��u�!�5PX�|A~�0��sC�& � �����2��}d��ppO�h���շ,�R���^'���^f�UmкG7B��s�3r�E�/��5s4�FL�����?b�s������)Ʉ(���En�˰ќEy����/�mؓ�(�Lż���