XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/e���f�Dn��Y�B�\A\W��jV���lN�%ë��hC�Ǟ2{ۦ�x�5��{&�x��e	���Nj�7�E�Pd�Ǚ��^�����F����<O#�Z@���A�1��Jv����d��L����m�g�M̆^1ż���1F�F�kf�8AI�!%b�~�%���ki�j"ޏ�����d֖σ���4S+O�� �:ؗE����3��)3��C0|-8��a�#E��HXod�
����xaa�
�|s�<���IazMI��`�aVLV
VB۾����'TF�8��ۢc(Mu�����y���}#�����g���zUU%ͧ �a����9ӧ�4;B���J�h�Z�j�L�N�$�g1�����r��Z븲�R�����Z��9Y����ey�w�-���V1����'�B�;��+FS�^@�2MҌ� �h���B�d�8�d��-�~>�ױVl����|�BN��EQ�O�c�plE�T��1�e�,B�6�(�|L��0��O�y]����`���$$���)�%�����~��H��x�Ʊ [�Gq��w��z�+��ʌ����ҶX!����Aҽ�^f�9����N�通����v�n�2��X���p�a����s�p�+��|�-%�|�g�qVO�����]tlj) -��`{�v��m������5E����ֹZm��eY:�Lr�L'\�i.aG��Y6��Pi��B٦�������jUt�	���Y�Tr XlxVHYEB    56d2    12a0�'R]�8�C*oU��ږY��t��u?'���k����=����Ճ�D�� 5R���\����K�\�$��2R�6�t$7��Qs � �$�Z^�d���0�4��)x��j�B=ԍ+*d����
�d%�^2�2�y�
%m�g��k���|���J�w_�x���[��b*����!B ���sJ,�	�ͫyUJ�e|,��D�����'�}��f�������^�L��'A�ɏiŎ�f;T��?9�W-��%��~y��	�0H����
K2�~m��(�aך�����@r���� G��B�b��X���׍����5�[�&Q��[ϲ���;f���Ţ�+���r(R�wA�.-�|nθ02� AKI� -l� �7��"���>"_VC�|�i��;k�歹:V�	bʣe`)�{��}P}eFo"h�g����/!|�K���σ��pZY�̕T��ݘ�2�h��d�W���F���o��r-�[H����@}L�Hj�l	Y��RvHpL�/0|�N������8�Xv�ܟX���@!����"�����s�_�^_���K��!!Jc��,!���ˠB�q�������CY�����*��ǭҺ83��Ͻt���%��f�E�������fZ�����a��4�q]�@��.�**�Q���Lw?1\����ipl��IﱿT�Sv�bgJ�yRxf3�E [�O/�J�!�)x.�f2e�t�:�aX�Ӯ�����gb��̥��x�~�C|�Uh5�VihP�0i��+�z��+/�$S�G�2�n�4-���nO�>j\���}0��d��JdP]�u�T��S��7R���X����dFӷ�ZE�I�5S��n5\N���Ϗ�z-n�|��Bܕ�氶�-��Nw�F�Mp���!#gݫ�TI�\�V\v�TD���`�e�o�0��rF��CPB�[FQ��&�Z/���D��&����Y�;iz�o�m��_��VyU)�&��'���]c��o~���L�20-�g���'�4,#K�/�b|�9�nE�*s�����~�4%�3d� �U�Ϸ����r;.��-���xu�	�0�?Sۥ_�A��d�i ��o�@C?k���.�f}7��.���,f!Pb}��Yl�t��6I��	̪���H��Bʅ�����~qH�es��c�q\��0��!�bVs��ݜ	X�f:�ZK����;N�Q�RXz\1S�z�6�O�bݶ���ϛ��r�iƇV��z��A�Ģ�m��Cr���Ϳ~,��������HC�55��-0PS��
�';%��M��sa��D��-Ng�FE`�M����e7���I�W��ɢ5��N$��]y-#�/ϐC�J����Z� |p�e��'1��N��3��[�Y�*0�Հ�Pu;m|s wR,��I�<��z����[���EWN�S&^`ᤎ�F����y�y�WA�+ϡp�(H�1�sb	$�m��R��]���H�~ꈍ��/�<���Mq���_�>*��䯖j��oMu������s�BNͣ�:'2r�F��:z�[ԅB�N�DK���}?�(�W�N(F���D��5(I`��j--�qdL�e�����x6_�g��wCy��g?CM䚈�U��+�p:����r"b��8e�a�n���O������9��v��{���I`�Ԁ���>��&��("�--���ܠn�ul�v��]w�n�Y,#�%sk�������0$�?�3�8\~(1h�q%��Չl���5@��\!�ت���S�aB���IY+��e
>�^������zS�~�+H���?Bф�����>o�V��ɷ[��xbc�ٕ`��`����t���f�1_l�-�a�ו�ac��=�-3�v�����፺����d�[n��s��E"ú�_6����<��,w���V�e�l�Լ�����H�7������d�U i~Zͽ�5�y���2��-���	p�tL.�-�& 3��C_���j�Z��9��~���TRV�J:E\G�5�e+��!�]�*QC|"-Gt�B�ز��bT���N��Wa
-B�4��+ۃc9JFd1xM�N@���f�����%�U�9s��-(^g���;����_�V6����v15Y�۠�4pWM��_,8F���Xތ�4�����Ȯ<@�ޟS���4h�� �Kj�^퐍v����o����]*�fly�!Eao�\,�kv]L?P7�)�F��r�I��Yp�:|�y���3bZWKK$��7O�_��s<Mr��ûJ��;��uaԞ�צ��z�$M��J�7�X��U��H*�i4	��T&��IK]6YGt"�P4�z!���L���pC,���I7ǁ�b`��F�C4���Y �HA4�M���=�On>[_����e�(��;Se��vF��%��f�;ԋ�%�z�Ug)��^a������� ����:.:�����6�����4�B�Q3i� 4��,�|��x^�ݜ����#�=m�h,G�ڕ�w�M��5��Lq���0yռ���~R�F��&����	⪕��R�&w�:���l=�e�IjL*+���� �4o��F�׆+��r�#Q6��7f׾&�5����u��M�n�0�ˡ����Y����$qX�� К] 9���Wp�3��:��+��ov�5���|�	�!����A�`)*͇o�x�~:{���wc�ډk}�=�˞7)�0X>�7$cE�gH~֭�_�F^pՔJS*V�!Ѕf$���
����!�"W���U/~h6��oo����F��<��Lٔ �@�XP<H]� �槪rm��`����[T^}�vY��6��?'Z��1��x�����	@��<��`�Nw��1�C)"�F�8p�����������~d(�{Oy�%�Ŭ1�E�7N�^�����5��㫼C��tcг�ư}?Mx��I�Un�����s����p��d���@�/�¢�c0�Z���{0~d�'S/Q�KA� ��;=|��s�4J��m�is���C
9U,_���t�	����78��޺�~�P���I�.���.�>t��y�h�(�-:ud�A�b�O!��/��a}.@1�)N�`�*����'Κ,3�#ݫ��	�${rD�m�����֍=�&����7��ѻV�v�a���R�w�K��nn���C�����<v�<b٥=��"��hq7k>��1����Z��HM[Ӽ�V#Nl����a0�r�+��-n������uؿ����*$�Ŵw`J�)�]���������M����^�f4vjD��ޣ弩�}�E�s��d�\�h�Ӝv������̄��Sᯉ�v����ԛ�GD(+wF�Օ��p] J_xv	�>8/�����s 0s'M �������;O%���5C����XH�����хRq���A��#��2��WSm��� ������!�x��������8�]��I�T$���+��DY�z��u����{����M�U{=�Wm���Pu[��?���W��nv'����8*���X[wU9���/�r^���.Ǭ`n�
��V��r�W�>*�*�����|���ߴ�y��3��{��#>�W<�\g���Kx�TgNkF��NHn����\հ�8t�H�R;�� ���2d8�*�M�dz�J����!����f�������ѧ�A[�%����ou/�����|��k�hr���a�4[b�7ϑ0�ݪ�p6$,�t��o�RRU��Gi�x����UƩ@LSq?@ec�l��?�7�'�����/�	i��,��� ḭ�AO�/�*�F��̜A�0������&�g���u&��-�uO8f���F�ꢾ�F��v����W�f�o���ؾ>����0Ӯ;jǄ ���{S/�_��>ƛ��v��=�lӌ^N,a�Cn�q����P>�3���	�]�[�6-�@ߧ�?-�� u<�n�r�� $9�f�-gy� _Ϟ�N;+�iˇ^b1�G/���|ϩ���������v��^���.5
ܱe�P?sc�H���S v��q��A0�\-�ߩ� �&�'#:�p
���,!4�h�����>5Y��Qf���i�~��}߻�K���+�1�[�����z�S����=Tҷx�ԡ|kfB{hvX���mA~4���ga�iB#�NH�K���۫��y����9��V��ɏ9]�\���=�f���\�ēi0'�W٧�R�����Y"�V<fT.����a'����np`�9֮/>�]+ey䊙EKR�����<݋�
�r��l���k�{�7伣JS9$�0�s[=c�b��{O<���}�����Vz�.W�k&�Md1���ו��i�z����B�o�![,��GS�n��>M�#"�TQ��L�?�Y��Nv,w=ְ��z��qG�k����8��6]9�Pk�7�e���[����$[L�%����S�:!����d�g�Z�f����,ŗ` ���� w"t���&%q�9����)b�e����0�������Y�H���Y�ˁ"oy�bX|dO%�&P�2:�B{����$�&����>�.����T9 V��j��mx_+�h����!f��v�IO$W��<k�����8�D��ٰjK]�w�aw4��z���d�+��-�[_��O]r�e͉�jE�'��$qk��A�Ok�?�