XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����TM�ƹ�q�����1d���.��`8���;Ԗ]7(�[E�J1F�m�Ñ�B���؊<kp��E����ִ�G�]U6�5K���Aʰ|�К��ۣ����"֔8/��#!�:���(x��煡i&� ����w���[U�X��s����)�2�"�O��4��F���fb)���n=�<eÄF�(�L��G��+~I����P44�B���-���.~�1%��&���z��絅!�����/�Rb�ֱ`���xr��L�Yù�=R;�D1�o�jS>�_͹���� 􆊄U��������R��w��J{��:2QB�c�r�rq?��;��]bn뮜��=f�b��z�l��/�	�Dr9�g��m6v�� h���2RZ`ѝ�[ԓ�p6j�����AU���N��Vvŵ)F)�['ʫV����P�2J6�j���-�$3�G��'[��J�߲�s9 8�^�T�/-'����[%�3�c�����]�4I��9��\�J�w���JI�R\ C{!"?��H�b6_�lE��,e�i�JNI�������=��AL�̏W��G&V)����rǓ�|�#�x�j���mJq@�z�M�LE�~ڸ/�v>'�f�.����P�r(n6��<�P:w�۩Y9�GE���]�MU��C��F���&��-a�4�/����
I�"��죩|�rc�:�[&,��$+ÿe�,�"'l7ރ�`�0?�n��H8;��lW��t3�J�tXlxVHYEB    33bd     c90��p�����_�h*��t͋ƨ@ܽ���#�TWj�B�C�}���_;��1.��[�"�%�Z�#�Q`�
i�h6r9j�VW� �D@x�yr#�'6�aP+B�N/�Lb<��zО�L��r���M��ť'�f�s�/w���I���ܭ�4������>���e�T��Ïͦ�-u��-���m�^k��g�,Q�����b�8us/%�ˑ���[�9o����U�,�@��ܿ��r	6g����$����>��i��zŤK������F��AQ���.��*"|�'W��N�`�����5���k���n��޽d0Z��)��}3� 3N�ЄP*�=�$5鿶Woֲڦ�I~Q���R��"�尼'n�E�SZ�C�f�D���R���5��j�X6���E�8M/�˱s��8�)x�����b���n��<dpK�X:x�d�0v��8A��$4Q��
�[�V�}�����֘���O$�͑���Ѝ<���'�0Q�_�G�r����z�L�2r�S!��5�>���,cޠ���~�q�U=�����Ʌ)��Ю�|%!d�Ԑ,����g}B��K'&��[���+�LW����X������5>�}ᶓ�70ݦP�dD�l�
&�{�������#���9goE�P���>�$v�΋֕S�����>/�θ��B��h�`���y������D�m����^�����BO_���)����^̠���r��R���_���ͅ��~�r;Ϟ��i�N�����.& ����6���<�����Y�RN���q�P�� P6w�AYg�%yᄴ$c���i��',K���QU��K%�r䧣O��E�2jQRD! u�!���z��~^�c��l����p����r�7���
�x(��\�+5n�3Ы���؈سQ�,�� �]�ʅMf���쳀��]Vo��tq�jη�c����1&yySJ��*��(��~6yuL��&� /���s��_*�C��f��Q��s������Qz�pE˝ZMD#�}-li1}d�1���9�G�̩��@ ���]���Sp��^�?4�,���Wd4����I+"�+��:�H�M�A� ��/��v����V�z�� ǟ2kxbk�R(ۗr������/[�j�t3�,>�xo"q���B�ߠt��^���j�#)K�Xo���r��c,HGrs<b��{8�	ƍ��V@0�CCŅ���z5c���m��n2��y'��<�j����}P;9��I{ʅ>6L�ǭ3H�� ����n\�E'z{�����3�vQOV�U1�{t���41m���wAڴ�^f)F��]3�����u*��L��BR�<��c!I;��71���&bp��+A�S��s��.q]
'mVܫEi�L5*�Œ���Оk8������^�눡��枭����U���0��EG�\h�9�E�♤1����oa�A�[o6���9�L{��E��j�DwB��,7	s�+�i��,��Yb��@&�|R
�J��D �����8�*��%O.��[�X��4�=LM�Vc`*��*�y	�`�5<�r	�oD`�ܻH3�;{��'	P�d��i�x�\f�HӾ�Q�Ɲ;��"[Y�Xz��l��6�NyTιڵ�`��GX���d��ZOdLXs���˲��m �S��3]X�P٢=��W�ů�O MM�m-��M>i�ě�y���͋�w]��m��1����sha�+�i�"i�c��(K�o�ć�
��ܽ��T_9�)BZG�Œ�k��0�*��D���cP]�FE'	�ǔ��|A	t���h�;BF��|zk��W߯��ۿ�ٕ�4�#�c��t�� �f<��'�9��
,����r6�5�Or���.�>�õ��0q�>���b���&�����(9�'3����id[V����[{A~9SƲ�(I�Y�p��[M�&��z��|<h��W�l/����7'��NAVg�ʍC�>�Y��O+�L�"y����t���v�ܿ�+���9?R(]��b�d#q����՛x�<����ޝ�R�U�!>��o�v�fAq����[��˱8��j���@����i��̀����4[7���x$�t�G�W	^Ł욺���`S{����|a+�`::Ip��˳�N;.h౸�8�Y�����~�K�g�8U����D�6�D�D�h�Y+�-��m[q
�����~��Wy��2b_��p���o�(�)�8WZ�v=��pQ�_bn��TQ�A��Ӫ�b��3����蚴y�ᄪth��B/\��������^�k���*5̀E*g�g]X	�{��=7�q<��X��~VZUt���Q�Z>��lt*<���Ă���q*u4���ߣ��Ӭ&�A�-��E-���ST@�҅��Ϫ>�v��:B�.siZUg�X�� k��BZ�7����&��0r�(����	n=�L�K]WOj��.2�zխ�܌*Yp������{�@���-G?�Q!�2G,��"�TOJ�����U��Ec�gG���S�"X�`WBA��,��<,J�-tN���7�M=�r�4}�Ji�G�1�=ۄ����������p�YR�����f�NO�X��z�B}hCD;]��H��"����s�\)G4���zQم�.�i���.ř�O���>�40,۞G):�I����|OC��T0�R^��44��`���,b#�Rq��ȺS���{J@O���pS&�+�nqYH@���6���c� )�C���W�,�u
�� �3��R��V1uz�E�k5��}=�)��H��]b|�N��	`���ZT����
���	r+o� �f��"\�(;ķ�ԄS=���b	ou��糇�n���\�g���ξ+�N��M��M|�n�@y�C2���~ngT�Y����_{ys��,ȩU�T2�`����p#V�]��f�Nf�V˨w�����㳭���C�f`X�F�8�	��U����t��"IL�ܘ�IBr,!�ꭡr2�Ӽ����h����:,��e��׸ KQ�W�u]�S*Ѱl�;3�t��6I��VK��|��l�U�(�
|�lB��i��? �r+��#[�;3���	��s��w�����"U�3��g��&	���k� ����R J��ktg���K���d*3���xE�4P��9����Qm K&�R��l�8N