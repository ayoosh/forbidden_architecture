XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!��E����j��J��U͛���.MTP�j�E���VӒ�J�h�:"�����o�\" 4)Ώ�v�kRܭ��k(��aR�tT���b�aY���YQ^���[W2#m�lh\h�Ew�����4����#b�>�}
�����)�d��>��B�#B-BY�9g��m{sS+��{��ow�x������C��<�Dwܞ*[��۔��8�q�m�4p$��=��U�==j�M�<Kt2��gǑk��_�B.'$r�׮(�i�_q�E���G}��㜒���_]8�	���ei�!V����[C$�?��Kb���8�{~�y)��E�v��d`9��,uEk�oBUI"����l����:�~�}�~�F�W�����Ӱ�������.ߵ+�<�����F00Iv��u�K�>��Xs�v���v?hf�s[6�>���V��(dm��:�����F7`>�!���T�$.����hu�i"���s�R���V�
�O(��^�g�d�C��$��r���<!�\��J��iG��i�~��w,��l�\�0�:N�=20�:�CG쀬�N�֞Y��c�ū]S.�?�g,(/Ƌ|�>�[O"����K!{�83(\J.ح ;9U�1�zͬk��l��z�g~��Sh&�R�����<�butK</j�� ��n��* Pe>�p�cIu�z�aE���$���\ϫ�^��4��E9n�o�::;6��t�|�&rȾa�LIO�ڤ�"XlxVHYEB    4089     e40US�u�
7ץN]<�#��僢dd�OZV�.�`��`����1D�)u2��G�������A��J�Y�L|r��q��?4���	�4kA�x �Erߟv7���F����L���j5R����r��L�ԻO���(#�˴·�9��W��h�,�C'$ă�C���z���5�6&�z�2�)�Ϭ�}��6(����U��@���R����mD��/!�H��~Jo�'�i胋_�V/�wՍF.(���pl���4}��0��:\9'U�_n�RW����%�O=��Q�^���o�đ�c�X���9 >Ai�i'�d�I*	g��aV���n�%�oi��d�4�#țG���l�ԁ�JW��&���|�ݲ/zLb�BC�:�����'=���%1��.-�D�����hܪ��ݘ^�7n��00�7Aw��04�{���D�	�檜�Z��_~߬�_2��,(wv�g[��P���9���A��0U��6:�$mEL*;�-k2]�z��H�绦`�� l�f;��cѹ�ٲόK{�i�9���U_��T6�l/u�^����Z�3i~�H�:O���B���ʅ�W!�ǯ�Ӧ�(�b�̺mؔɚ�<Aue�. ~K����k(O%�/X�n��`�涗�ўQ=
�����Gtk��Ty�-?�N��
�'�Ý���B�#�k��F�y�h�r�k�v;�#�f� ��/D��i�L�"\Z���t*\lq�0��5�>S@Γ#U���4S�G�{�o�����]wD��Rjkv���}�@�U���'5kx��2��UU$<��:r<?�3��q�.�U�8��<4b�4��[���	ɝq#�L�9�%�T�d�2�v#Wf�B�f��R�뉐i��i����i<_&�p�u�s!:�!�L����L��*6$�2V��Jl?A�?F�3�t�X�w�ʂ	a �`���9q�A"@�k-_0�Q�Ytd�pu�?�4m��ݥ�����|I��TV�R"x,��_%���j�@ Y���-F,LhKnt��	of�֞�r% �o����be���w���Q�A��J���$ς���^Q��-nF�j��v���%��Cھx��ulk�t��]��\!��x�b�d8hzJK�Ѕ����.Y}m�J�{6^ �3:P(���}��X�=��g�M�Q��h#ca[��������Ct=�݈0�%������\��T��>d���M;�_�����P��a��U[΅�@a��#�yW�:N㜤S4;͍�T�2D
����)�x�ypa
�����w Q��!>r}tZ3�c�#�$Bg��^�^Z��:��^(��7�wZA�E@Rq@My�a����"�w�9�뉳�XOW��d��N5x�eD�:׭�Lq�4
xr�19o'�"{f�e��)�W�_��a�ex=���%h��LP=��+�w<� �`>��'S���^,:���~�ۀ��/�;<+	LV�텱f��(��ۥw~؟Y�[��*��7����]���qy�x�,�Qˎ~�l}D�%��^�l7h����j�EIh�6JU�Ym�*o���/��eik��^���(m���Ǥ��DIzQ���@J�<�R^�ь�~k=���L�z4 ��MT��,-+a:hɮ��h��9�{E��!�S�C�,�	XҺ�~�@l���v.���f��U:�p+�.7��B�����o�������
��ܱ�5��D;���OJ�ַ�$���ʋ�+��Ȉ�&�H�3Y����I�Y��k��d�1E:�K�����d?�U���ܷ�wWQj�v���.���L�:G��bFw�ֺ�S�c��x6jae]��7�Hޚ?�"������߾y�g�J���'�a`��w*��Hќ�-�����,�`�_���Mh�e|�4�V���i�:���j6Z�����Yn�k�� 4�pF_o$�%���Ǥ�/�UPo�L�����4��<*p��o;љ�Y`�Z1�h�n����_��e�(xH޿�yO�z�p0򳱗�O����f$��T��@�r˧d�>Y��U�P���B-�Ƴp�l�zΏ��ed�����&�I�m��p�}���N�Oǡ��k7{�Ͳ@=�����K�<�[fj�m�QI�{`Qt0f޲� =�.6Ò7�I��Rp��w s��L���챯�U��sj=>֛�/����!���f��(*�'.�S�ҟ\�4�t� �f�j\+[�(��!� F�w�-=?FAqP`���%�31[@ S�4�y"��&�@3:Ē����K&��"��B\�`n*tx\�^�:a����e��U��a"�>�0��2I�	��	9^��v)̇���\U��^*N�nM�9����=hܔ�j��A�i���x���g�����aMb�>�s��_��:��C�s�2�߬*�TI�6إY<(:����ш�j�)��G�'�=����`�,	�����yR��^�Y,�I�oˤ �f�`���k��-8|��@3��:Z�����4���V�F2䷹I|��R��w�m� 46��8��6�QO��|8v�>�>��ZibI�I�����<�
����n?-#��/���&`NI����	p�Ɉ~����8�`���GKV��Bv��l�I�"�Z���2iO������Y����4�$��Tί[f�z��u�
��Ma�\�|�0=5��Ka뻷a��1��р,�e��
�XWr������Aa�����vD/��'Pdů��;2D�m��ǉZЮ�):�J}�] Ŭg��'�UO ��jB�eJ��^`�Z}��
�|�{�z�b�8��=��%ZwMJX�+eA͠�%r�?���Dpd!~�����=[p)ؒV�0? ��������-ўQ]�Te���u9����4����������"&�喘�);ι8K߂����Ky�:��_ƹ86���.h��j�s-��u
�}�S���UY�Yp�̨Z�Ž81���'��ٞ\���?�'~Br���ݰ\�"4E��D�������H~ձ�^����\P��xT��](�o��kI��SA��W�N�������[��<F�"%D/NZ�6rڠ8��oÜĒ�1J�|�F�C�c�g��a)�fv�D#�{�Yi�b+7-V"7m��#~K�Ե�-uR��:n]� Gw�&���<�.�`*���Q��X�>f?y�%z�3+#2�D.����#���rH?o��U%jS���`f�fL�%��$�3����L�+8jz���n+Î;76d��Y�5���4q�]S��Cn_���#~�h�}���w.��,����UN�t]u��$���Ev�������u9����X50uw���}'�?	q���E-�պ��wY��}�C��  p�ȫ�4��� @Q�X�h�x�V�*�����{2���4���Ѩ�B�p�d����e��4���ar��=�f�){:'.S+1��g��wU	V���C��L���4@1Ɉ5	f�ZlR'�N٫G��o��m��F�3�*��a��g�@�\�������H�ž�:�~w:��%��@�n%sG