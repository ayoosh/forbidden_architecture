XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����A
N4q	̴E�<�!u��P���ڠ�\+����+z\_I:��x�v�B�8,&{ʙ���4����J����c�p/1� #N�a�=?S�t�a�!$�fx�w��W5�.u��C��,�PG:��>Y��5���oF���ʀ���8HO��qW����O���R��-�@��MF����	�-���X!-�YV� |�&�Ή3]S�c�{��tV?��	y�e;�,���M�16O�@�r�'/�-�Ú��ڇ���PsR����A@H�D0��(
0������O�/���b�D�VA�ڞH���Lm%Sː�z�q�*a6��f�s�A'z��ӚxQX:���Ft&(QY�8<���}����G�bI���BF����km��B�lZ�]5��{z=.a:��!�)����UF�b�ǧ����\�� ߶iC�.v�zȁ��K>��ɑ\�-I�k��W�p�	�Mmj\^|�#f�`~pC,����FM	G3r %~~.�v�`.���|+��)冗O�Z����U��Iܡ��|����;�}��h���V1zQ��Ig��[���kc���u�i����7�s��D�}��M:a��4����֣ϼĘ6!����f<�ڶ�I���rbG�^2 V�J�4��R�V�z���خ�(��5.yh���#�Q�E'���Q���#�0�k�\���X+^~^��@��Üc��4S��c����w��̍���af�=��ע0�����lTXlxVHYEB    8e66    1830�s[��]$�P��{:'���- sw3ї�7��w�A9�F~RI��z@�v��	�5�6�:��0�De��^d�e�A'�I�\ِ�E�-����Q���N8���	�KTm~�/^=�&VƢ�ك(k[5�]Ҵu;��mj!��Ky�u����?�5LԠ�P���$����W�R��`��*A�Ya�����61MZ��E+��vwd �$h�3�7� ^]G�*����.�p>����֞=��L�)B���:ͨ�qx�`��cL�o�����|��0!؀�"�]�k.����/�A|JE4"�c��.��EM��X�+
&`�`+�Y�Iϫ�.؇^:�ť^�AǍ }̱xf�� ���K��_M~nBo�q[!v�W����}n��&i��0�S<�A��nIRّi��3���TÞ�.$�yyt�7�6�����
m��9�W��G�qK�R�ns�2��֧%~En����Kiw�R���Vxbg���EGp��V��1>gZL�\ԙ&��?����W��
TQR� �oc"�N��O|�8�	]�X�`nJ��^E_���gf�EŶ$p�ay��G���JW7a��BI�u���������LF<9��]��4wiN�⫕M�2����� iv+�f�K�
�>�Y�?��5&'�O4�&�ݱ(�[�&J^�*�_&���o��:�5Ir -�Ȋ뛯�w��8�;E��:�y����n��g����	U �w��F�0�ǸE_���}��=̑��_�:������ �ˬ@��4�|h:��1�����x��qu����R�hV��� У��5�S�;��zY�c�2�j@����F�Npe�R�����<~
�f���T!|�	v�w�D� s����LM���Q7��}#�G���q�7�|t�Mc/�1���+�/��M�6w�ݞT�NMC�+�y�ȞPNJ7�?��[���oWac�u�qv�h���x88 ��&?�t��P�h�W�����i��8�O VA<�wD����I�AH��t=�	�i�/��V���fnG���fq1��,����h�_��z���]&4��Lx\�j�o�_�4��s��v��s,���R�z@�Uh��f�W����C���s�U�E7��}�ΔA��w��
CZ.s���qe��4?8F��$NI����u��D��,5Bk�kX�A�b?�/dB��GZ��i�8�լ��U��Јh���#0{\�J#LU�F�f�R �<qe��m]9�e�w�z���b��%����t��E��������yAs^�K���M�j��B�x2�
�����%��mw�(�^��%��7LW=����11��0��|��'7�]�ld~KY��^���Scw�?�u+�F;'�N�(Vܒ��̸Us6`�� e�ĠZ탔��N̎țI�5�O�}E��k�_��w��}�~����(^�����;6`Xu5T=dQ���/Q��8����s�@|�8\��K�uf>@	Ceo����$�?ў�����훧@*
�~����G�I���:`��� �����>��˿���!ٜ����$8���d~Jb3�X 4B��w�e�7��a9v�eȵ�j����@�s}��^ �q��/�*U�?.�>��"���f��Q�^s�Z}���ym�nx�Vv���V+�؎&���R�\��J�g%�v�����tA?������^�;�������y��{ɆNہ޾86:�iu�}�j�"/7�^Y�%�j�P�+YH��� �v=,�kg`=�~�pOts^}\��0$7�=�읞1Z�dZdno�D��+њ��ęol���,Y0c1�FK"�3D3)-���9Lk������e��%��`��*���)R��vF��W�7�U	����妣���,i���ݬX~)Yhϭ�T����L����֕�-�}�m#;�v�@���i֕�V���'���K:�x����P�~�X����@ш]����bR<˸%���V�E^�`�huAK��Jϧ��t�������0���N����/ד%�<̊�o�w����oe��	�`�qqh]���A^=ڳ�N:F~8Q��bbtN}����2OOg�l�Z��M嗅쪓}�@_��'*Om�/��s���6�ǝ�0qZ�ԘHCF�������l*�豯UO1S$,#���E|
�K0�U,����B�IF�G;r�6��}M7�\���-h��8Յ��% ]�ӂ��PU>��9����ē-%���(�p��G�C��4t��3�l�B���_0�iR���4ߙ]q�Ů��s��A��*&9�g�����-tn�fPCT�{�b /�X�����q�i r���.����6���{ a�������A�����]rb�����Uu��=_���x�M���cb*g���!�8fąѕ��v��2�6��XW���c)|��#�N������-7f��M���)l0��n|��CR]鍝�N<[��~�Y��έ�z�l�^Q���z����RH��@u�.�ٗ�����U2��n/��]R��� ]P��2��ϭf�K�i�Tc�������/%.�	<������>^�~ݧT��rN���]a�c��=�����12��,7���°���>lq���p��L�$B��c�/����3x��i�sj"��L�Vs�)L��QyĪ������^�ļ���D)�PY�#�7�L{�w�9�1Z�n�y��tAw�l�t8y���}��%L�ۂ����9 ��5o<�מ�Ǖ�f,���`���w@�^��-�t�#Ѯ����xD
t���-��@a�,�y��y>�Y8�@�\hl#A�'6D]b(�؛���~�]��C��0�$�-�p�r�Z ���r���ό5ʖQH�`U�<�. !���ip���۪e(� �Q��uU�� �<��WR��ʚ��ȍ�O�<Gj���*�`<E�f��;�.�UM�2ۀ�-�������X��*~���3X�
��˲�O/���]#Yk���U8 ���TR)�s��w�ULw�U��jǞ4T������ĭ�ŏa� D꺍ό�u)��$6��@L�mG��ܛ�O�z
ғ޹�N�ӵ:�x�����utnY��;:�{��ӭB�^;�Y',�t������%G��V {�r��l�$���]�A�0՗�g{�l���a����Y}{r��i0��Ϧq!�{ ז�9�<��t@c˹H�./M'��54/���h��G����E��L+�T)�˄�o�ͬA��q�GyN�6�/�;`���������Q��	�'%�,��5�1_E�`��>�}A RL@D�i��e!%#�u���p�\N���6�Bi�C��q�L�\��]E+��zYc!����o���)
'�8&����=�@��r��`y4���"�_Qx��ތ��\oONHl�<�S��Q/'Ǩ�Oz���9xWFY�&��^[��U���P+����V�5CUr�Ax�?]�=q��|�����K�ẕ���T��2W����C��Ӌ��+藍 �G�ݯ�NY�+C]f�+|�6�>�r�M� ʈ����a�փd �Q=��m����kz6�^�}�QȠ<*���?�W E���E�&7]�|��VC��	�~#Jd����q�*�(Rf.�Y�b�}˧����)�cR�(>o񀊦����9� ��7�L�p�+�B��t A�~;p������nU>�}�D-�Б�#�ӈ�ѠH������7�-�"�Mq��I~w�%~��#d�b�]�h~�ޒ��eX_��etP�Bd��p�I����n7%�wE�W؀��gf:�)�Έ8du��8Z$�9�i��Jة� |G��%�����-\J��ч�P�un+;PnZ��~�]ާT>��,�a���g�C��l 
�iYE�� 1EX���3 F�4�FF��%C�F?
 #�X��S�����ζ�CW�	�@�*�ai�T��9l��)���](5�SB7���8M�X���]@�t��5$(Zq{;Y��h�~����>��g�a�[oM������6�"���pZ�:]��E���E-0�	���p�9�y�o��z�}�u��Ѫp}6�œ��-����} 7�0"�yh��� �+�5����.�u���x䗔�38�N'��Yt��^����nd>#��r��B�{�5k�U7uRQ����]nbY����ˁ\VN�҃0���%W�M��➹}��Y\<sڕ�+a[R����՚= ���l���ȏiV�A�*H;���f��h�@j!��^�)���;� ��
��q4���U�!�<.)r!�����q�[1:N��F�gtƊA��H��i����H�Ji/y��A�G4�JQ	@��D����:�]©�r���\�-�vZ����� &c�:�!�Y}pML+�"����1��S�?ǜNt�숬�y�X�-�X���vf�p��G�Ws���҄,�Spys�=l���a�B��5�ّ8U���o�Hlv������;�l�k��Kg�3��H)������v<��r$ia�n�6��{��l�T�%N�R��.y��ؙ�� tp<�B�Q��B)�>�R�K�����!`W��+}�@<�q��ݤ�X����B2`�_x��n}�����A��D��~Ih�8<ם� ����b��Fӯ2aK��F�S��m!0N)V�XAĸ�|*5i$̡Ä�"���AZ<P-�ɳ��TH�% ��n��>m+�(�gzDj�[cbDԥ�*��'�P�o]W��(�n֕�ɂ��<��,��jŰ4�2�b5��!�r�l�q�(�Dph�[䄍G	w�G��ES�QJ�u�
3�5�e�{Rϳ�<&u�V�:H�G�Z)X�UX�%��ňk�������s��B*п�>:���C�&����N3� ��!��Acz�l��a����M��;ǳ�_*��R�������up{	!�j�A�/�6�\�,���p#Jl����g�&�ݝ7�cCI�m}�`Wұ���~�51�6�-��&���;/=\���ߣ�x��)S�df�����6;E٦�g'T����+�o�V�\3��T���zW�*O>ۍ��R�z,
:�V�X�:���Vq=�~�>X��w��5%O/1�f;GC�Zb�~$@� /pt	q��{��z4��,�.� ���=�2���A̊C�3�kˣ����F�@�}h��[ޢ�CO�J�\ ����0Y��owzŚ����e�����ή�E[�N�F�:Urt�.6��ȗ�o�<�\c�`��s��{�(}iW��K���`U:�H�'��1}��~i�Q��ɭҎ���vH1�6������C
_�@��ř1vV�d���}EΎ��7���/�q�����ή`ySeĞ�*iʎ��B���(ť(���c�/4ڃ����4�����GC[\*�.�K^���1}S���P��j��C�%)�7��$Gw���tm��s��лS���Z�đx���ʊ�4�g���d=ⶦ���I6��#�Z�_����( �ce���kǜO�RΑ
��{��zj�;n��)���aLZ�ƳDV
l��w��(mP�8m!��xqlr��ĴoՔ�B� <�S跩	���zP�t��Ϯ8����u��ˮ���7�3$S͕h�V~�>�78��C"'`� j�)ǘ׬�MV���OBOl
p�����`'&5o���,���ro8�~��|��K�	'bl���� =O����?�ق�]����q��,��U&54��W�q"�d�� 9�auY>�=�ʞ}8엲_m�oVo�M~���ڜ�R]F%REO�8o�·V����a�9�Zת)>���q��O,�����Iڵ�ǣg#�P^&TK 1��B�jm���չ�N�P-�a�YS���������g��wtER�-����>��D���k�� Ϋ��B�\_�蝈�㽯��YH��A.�Uzs�޲.��8G"y,����ҭR�F�A6\�_�TD�3�\�o2W�������62��e,A�xo��+C
��L��