XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H��6�����.��Uѳ�!�(�Ȁ��v��h�/�'7� �QB&'����1*z&jCy����6��
=j�B�d����V�hv����YݕQݗ��ϊ�'�Y�d�_��s'^?����Lk��a�M�Y]D�6��>x�Y8�S�_��`��p���Dmic+������K��9c���ZG31z�?F˴U�ƦV���Yp��}���2����]\>U�/Qb�{dU�S'7��>�
*�af��/����7�P� 7����=����W~�L�mV�=��QL�(6r�#<Ox1�m��fӀ\��;���$��v�(�1�|H�Ԭ ��|/*	d�״,�^��7{�N��Y��630Т锔�o�N���f��t��Bـ���J��+�9�(�Qv%M�f��%k
ջƮ���2��Q���/6~���}�7$K ���:��5n/���V(�:`���>�v�B�yU|�Y`Gg�^��,��6����n���[�2�V��}�"B�U�F��N�6|��^�;y~�⻼Dhek#c���	-�RN�L�,��+p{v���s0D�z�>8�����1	�&1��p�ޚ��L��dr�j�z�|�	�l
g��.��	��/� �hp�:
�L(�܉��g��z�=���&�mk����c��H��轱�q5*��2����5�
���3'�@i�tn^Ǫ�An��<f@BI�b�$���p���ǀ%
<�H(�ՙ@�����ߞ��u�zbdT�@�8��ߵ�,��XlxVHYEB    fa00    2470c��?���MS@���kI�h�S��=��f����:[H�)q��\�K�Z
qp�q��k%�JAϺ�a�i7�t��9����[�J�!�Ar�5º��1�Y	��r��l�Ѐ����yX,�N.��D��d;�W"���kt�O��ր���O��U��%�u�s�/l��Ѫ���[�_{\
����|O{���� ��u�Qhy�(Yd��|��~f�/y3��5�֒F�i~��9��6����:$�0�Qmޤn�J����9���əl�e�4���ÔaН���ж�IaB=�1;_���F��;)4��K
�jΟI5����|�ɷ�J�4|Ja�[�7�b���&S�������j��\ԗǷ����Ʋp1/�Ù��M	���v.�:�>i2�%�C�%�2�d�W����#����L/2uo����{&�K�U鴀�ͪ듘�O�e6o������3{��E�pGS4y]��?6���}�Ǿ�H��nv�]eچ���t�!9-��S�k����9a�eQ;&�#|�u��V^v��x��Y8�Ԋ��y�/��t{�G���vl��8ѕ�hN��f?�/7�nE�e&��W��oz�h��z�̩��� ÁQ��r �3C'�ò}�(�Aq zv�Y��&OV�$�mi>�|�;�ڰ��{�6$��#si���m�_��������u#�4�D3�{!^�������Y$۴t�K�.���Z(�g�/�������b���`[^����él�x���؜� ��Ѕٔ���{t�����SOC��r\���X):�j4AՉ)�.�c����/D�#q�m�2����ɤ�*b뽍��	��D	8T��>����@2%��|��5��ZPUZ�s��T�fXpq�
0���o���`Ew�b�T��-"��O�	}uN
���ؔː�ÿ���~���1����|d�7��x�ƪ5E`7^	w�{�p��Ce2������V$Ey��4�ޛtxZta��J���u��"Ԑ�`ƿ�@&H��HV�<ǔ���{�pO� ��΁E���[ӝ��~"/�;�MHX������9vN|�f3�\��E�}�;���U�P����$�ӱJ�x�>Y�N�d��ӥPaXU,_��AX2�R�p.i #Q)߱��E�3/o�Z݉���K�cP�%�7V�����Z�>2pu3�B�ڍK���H��`OƽjASw<Q�ֽR9�C��Z�8V�c�J-�$��]cӸܽf��Py(����K�:P�Χ��%�T.��p�>z��2�V� '��+lZ�i��]Vn���>��E���@6��'�ʶ��M�c�}��4	X��s��̲�w85t���W�(�#�c�E쒠�eԠ�
3͞�����i�8'�I.��nB�Ʉ�i��I��j"hyZ�Ӟ��3���n�a������	��q6�9>C5�]�恜|z�ڃ�u�����!�>�f�� �~ЮP��­+�'bQ��7��P���2��pp�ꂄ�së��v���;�\�7,��n�4�n�Q�2�"e���H!.=�sp*a0>�H��7��z��� 6��Y ]1�����cA,X�`�ͷ��W��{���2�p-��.���ފąd�Ŵ��r�4��.�����P�ЌF��5ro记:!䴥Y\{@��b�=/�ˁ�Ղ����h�7�@q��&}F�S��t�rV4,��۠qt�>�;l�6�t�:�[�JL#��H��]Oi��RT�m�X~�y�������	���,�>��9t�Y��K�?O"���c s˙ӳ<��m�B�Cv�R�;+䨍2u���ʇ�&xr�t�o����x�O0�$�`_�$�*�(־��	���T�m�z����*U�#e;��?�Y�w�.#%�4��gX0�'V���C��9��؄o��Ⱥ2/0��k�X�^����̧�j�e�R�B�Ap:A!��@�^�BX�f�q�H��`�_���{�3KGn>`}g���Z�.�C��`�e�(٪;�����2xx�P*��[R7S�8��d:wя�\#��٪`n�U0S�-l��y�I�e`)�*���^~S��-%�w�|��pǤWɰ��Zr��[���)�:+���A�o{�R� �J4]\��a^P��GJ!�.��~���[�	���q@t�ݮ9�qs�y5м4�����O���P�z.��l⢵R�^h�������Oe�*�NQ�;�s�D
��i�?��}�Q����TI庛9hȺF>N$ai����!(s������19�uNt���S�v}B4!�31��zfCj^����EO(�'�c��S����-�^1�Y����:��r�΋X���a����眩9'<?��������zjJ�2􎈝Ԓ�7e�H�ȠJ%^YCCfV�/����׫b;�����EZ,���-Pe^�q�}�p����ͷ��p�ftqpj��M��A%X�z�����c��o��^���)ߎQ�5b%7gW|��]Pr����X!��`=�-b��ڡz�x�-ڴ�v;i�薒^�.���l1�m��9��_�j!���Ds���+cR׿��}���h6�;�%�ɜ������ ��O�c-'�Dʤ��ܝ�a��Q���h��}�N3\U�}>�	�����Y���L�F������0N�+����b%�.�V�U�%Ը�}܀�?����G`�8�3�9N���r-уm�1��:z����!<k�(]����z����yKe�e:C�T�'³����H׬ԎKR�'G�N�dH��1wB᧓<��r��?F��\�y�H��^��+.F]  wʮ ����N#��m�I����~z��癱�la�Ȳ ���`8<��b�������{���������	�B)�U^[��St݊�y��n�\�����~�~d�C�����g*2�T�r%��G�';>�;`B�f[-K���\S�8�D��VT��~�T����%	�p̿x�D�(0=�	��uAŒ0�y�-w�v��@�50�_�g�; �w�|�*d4He���%&z�k� r��7�:]�Z��MݻZ!:By��]����5�BLS�M��F
Z�O1l��g.�����:�e�l�s�:b�D��\�)���}4z���c��4���t6���a��X�R)�>{����YSsc��llIz1�'���t<�"	C��8�X�� ���=y��#�>j��,F��MW���rl%�c�����R���,�\j��ܸf;�V.Xh�m���A�m�.�S�����z�!tL����NM��3�[!n�>D�~9��:��Gv��r5�1�5PI\_�o<��cY����z��Ext�mmI�qȧ��l�}��U0�9Կ5"��g�R����>�Vr$�����Ν[q�݉���Ӡ�V�Z<U�0~����$�I�h��{BS7[�JK��s�iB�<ubD����$/jF�����&��M��M�BVFQ����D�`dL:H��޷(����d�Z��R.��WV<�P��!�>�{��Sj�9�F:�$B݂ T1r�;����H����-p߆�&61����o\����Ĕ��b�!�� H�g���۪�j9J/l�J���3��AR(�u���ᛊH5��F[s�v��P>�/Z�[4:�{ǔS�I\`�Ϸj`9w�е����*ՙ'��ՄE3�t�Ģ����D r���S[P+�jV�+LKO���wM&�Ǳ4悱����o��ۃ�Mq�m��`R�)B�M^Z�r��1�߰C�l�0�i|m�T-C$�uTg?���i&�m�Ҷ�_
ϵv�ä,<]p���b\����I߸!Qu��x��������`'"�����z�r�w��\j��{ޥ$c?5�9UkO��;���(��$�Ƞ�.��[��9,���q�1�d�D �ԑáB3sG�xR6!���)�4�-F4��k9de�^���4��:g�lV`q��u��iojw�ٝ��Z�`����;c�w�x�d!cV� jD���dю�
><�Gn�@�+�꺞�C��a�N:���\��vu�bk���,��Z>����i��f�I�үs��*Ƥ�1����5,M.�v�I���ę�@I������\��$s3�2�{VfB޼��:%���|ZY-<��=�ߪǽ8��U���kF6r:o�N%�3��� _�O<�$�m	@t����u��V=�n�
7¼�*����w!���4�+R/k�XX@����>3��$[_���e[�^;U����A˦�ȍuC��)4�u��R�A�����\�oW.�d�w�&�<*��&U]����b!I�A#�ݪz�&�����m�G~i�N�oR����>��͓4�5`���+��җ�y���&�'���%���T!m�Њ���c�.��$@-�0��i�L��L�����R�K#�]���]�| �k�p����˯f�i�V���'V�� A�����jԑ����{�ڼք�����_M�Z��A�'n�����[I4�O�0Ũ���:�c�̆�c�1Ւ]��\_�o�Ք���h;ɨ>�գ��gQ��B���d��c?�:OO�_<��*|m�(c��&-��_HJ��`H���jR�&��X]G��O��NU-)0ċ�}Nߎc2:Z����#�*���*�m5����t����'t�62�_�r��m���a�*y��Grv���@ᨰ�"���/������5��Aqp����i4)�9I�l5�f�����J��QN��!�N5̀Bk�o�s|�Lj�4��g�)\zLf��׬ŷ'࿸k��?gՍWu�,iT#����^�bG�����4��-@��ȸ����.�G=Y|QϠ���GJ���$f0>���"+�q���k�A~�(�m2���(�&ࢡl�c��+�v��o�=w���w�й�8rˋ��Ȓ	�9$״�y�$���[vM�#�q�����%�[o�5kLMT�9��'�jV���7��������$��L�IC������$�7��e���됌&h�����s�Ik>�h�ǫ�Q]�RʁʂV��C�<����h�����X�#%����M p�RLwA��6F�ɀ�AN�Sǜ�D��s�(��nU�fd��,��� [��埕��~�'�0�4�yG ��,�;����Oe�.H�*���#1���b!�v�҉٘��fy�	�ӭ�_�ZرR���~�f��^m��'JP���ڼ�i~���9�G���f�)-�Ӛ\B��.D�����b�9�7E�}�s4T�g�7C�O��w$��.<��>��ׇPr�J�rK����qB����e$-���9C(I�lo����V�5ǥ}u��7q��"
����ơ�k�V��V��9A�v�	xaG.�3�Z�񤈦{�Z�V��*����>��P�e+`�C2�ybZ"E��:ڸ?z��<�P�]�����<��#�N��;Y_\��R�O��]W!yD�`�����J�g~�(�{�@b�3K-;,�,�5+�*zQ��࿡��Tl5��m�xjD#Q$yC<�Rzr9���7��������A�A��xK�lK}���nx�n�'�7�1�_��t��B���c�c�ߩ���Ɗ��fZ!��(YL�t��3�l':mA�ߎ�H���^nw;fmxK֠u�rЊ���~oR�8*���&�.�Y�Y�� x���,��<T�z�\ln˔�"Y�ˋJ�Z��m,��]�F���i��lP%в6�>�	���RtY��y��k�jsm��E��;�z|_+�p�y�0�h����4>�r>�q~��w|��#�,ބ
N!��2���
���H��Υ�J+����3ፄwn`�j"�d��J��4��g~r��a.��� zP%��z�a�瑵_���ڲB݌�O�|���ūXYݔpV��Ѵ���B�.�G����Q� ��C�������R��scD�ζ�·��e=�r����p�j���=���>P#��� ~94�g�&�Fq\�3nƩC���	���VA�J+N�>w�	�Ӿab��a� ���v�Dҗ5����<�ǛL�g!�R ���3���]8�������9��խ������ZL*�{����\��?�U���z�uqFqQ:�B�����R��i���~`F;����6#Crm�B��n�͐U��I���K1E��#� ���w3M8SCϚo����3N�,�wo.��܅ɛ_O�S��5Ln�h $j��m�\B1��;V�iM�gWp�����1M:�J�!6����7���pYg\���zǸ��^`((|y�Be�{��1��b�a��\T���-]׽�/03mo4O��)U���M
���1�AC#M�<.W��7�m���r�5t�C3�, ��>��j)��R'__��b'6��X̠_ͥV7��N�)) !�G�G�̴T�B@F)����)������i��FK>	c��D�n|��X�n��s&zն__�8~1G��A�H�B����&� ���}88:C����.�Fu4�>�Y���/H��[���1wHk/x�����F-d䟅���3��>���~/�5�]<���LՂ�����Mz&![,L4,��=[�feX��%^b]�U�N��������<���Z�I�����3S�����\烈�Z; L_�x~Hf�7�����h�9����
�1�-��h-]Wu��Z:��S���o�BmϺ�X�h=�t�7���m�'���)$w�-����q�#��ag�[>�����1�qƥ��.u%fE p\�9ߑ���9+�1"Q��/�GZ���2�x�xݷoJ�F}���=�������ûى2������4�2�3g�d�@��d,�FK(�R�$
|�|�	pW����� g�ƭ~QB�c6M䀖�I�����z4�n�_0��e>�h9xok�.*ư��g���*r������9z�Hι�bzz���R�KH�U���naE�������J\��N���و6`g�̊J^�c���j$z��k]||iy��oZ���O�����ﮞv��KL�B�X�3r �����`.)1L��V���R0I�V�L�n#tM\%��ߴb��$Ȍ��]��O�q� !�޸r�9�~W0��)�~R)�\�20�gȚ�tp�!����_򞞞����b�eS�{�Ѯ�W�3��U�ӧ�cM�u�|�Ɖ�($�Ɋ�H��T�M�'\�[J���M�g�H'���\ K��2��2�����N�Ӡ�X!��8��ʜ{.Bx�F�%@�	�Yq���W��1
02O��Չ}(SĜx���A�2,J&��	��.Jd�DJ�7���C�&=����wC�۰�Ӻ1DdQZ�a���"��N��-�ϦIMR:\�ޭ^8a�:��*�Gs��Gu8�׺�Wܺ1hѲ�Zۏ�q� U+�=�ɿ�F)�# UR���[��Km��/S�E}�|�1�L�q��v���w�G�����SBJD}�8�8b�����Aې�/��Wjp�=~'W�ú�3����0I�G���P��mO��|����̞���v��?F:#�`�*P�܍h<,(�t";�3 O�����j��30�vϡ�ʀ^J e�M���W[��E��F<�[�Wl���Wm��#�OZ|%9��8[ޠ%�N�-��<��Z�}����q��sg�(��hdlV<rsܩ=�+=�U+�$��Ϙ>���[&�X� ���:�/H�4�Ȅ��c��.nޘ8�����@�:��F!��T@��
U���Q�����q�ů�0�~g¯΅	�t.t{�=���m�]��Q×QZ��d������Ҹ�Ad
8�:��߀�'xIN;��o�P����,��Dڔ��#q�ؽ@l���s7�u�ʣ����-�s����N�9N	p��T�骋z�m�z���f�ܶ=���L?�y�U�[c���$�Nm�\�B���+C��\�9�����)ʼV��!��A�u@�g�ށ"�vW�O�������f{-��K�7��J�L�b2�e��R���{tF׍�olnb�j趬�@����8���'f��i�1��2�/�}��$O��/UN��^���c������~��nǃ�����`���	���Rp)g��N�1:��7��T��dGP1'C�6��UV�+��Ԣ*hE��:��!ɉ;b����4��yY�?�H��Ewd)����.i>~c����De�5�R7�`Ti�+�LR��5�X�+���oz�=�e4�x����T�3D���6.=�!�)C�q�>Ts%)�>�[`0��H0�͸JS\/�#�K��p�ȧ6�a��r9�R��F)q��h����s9SX/q+3;��ʯ$�=�y�+u�ᜓT�у^Z5�e����\��~�9Q�؄�~���>�SY*�>���˃����^F��V.���\E�<��?d���z@���PP�q����j+�:��~y�؇��3
]���2��~�E�@��#�ֹ��kރ#����y3�s�g��)�SWA�#�#������)��8�؜��hQ�_���j�K�5o ����Mr�q�$"p;4���"%Ʉ<9x�۳���0�A����mʙ�L[��gq@��q��r�p� ���b�LL-h��5Zr�B,���X0:� �~�Yq8𞋱x5�*�v3M�/�;
���	��3�Ϟ�Q�вӬ����G��[!��1�5��t�L-]�3o�=sd��ݻA�㋆p*��/2�Jg���P/!�D�/h�B0��.�q���x��j���:�SDLRvu�n^xB�*l�ln�8�	�`ş�)�x����c���ɰ|�F�4�N!Xo����G��T��$oe��\��-a.�w�L�M�Uk�gؘ���ws�?��okʾ-�6kP�M���҉�Y|s�C��/��ȟ���|g��b�[>�c��Ab�֒Ǉ%�  Ŗ��~k�7�����>���.�����PN_�	�=L~B�J�<d��s9�zK��ʯ-k��.ˆ�,Z�?��e��[�+	قA�ld6O�UN��~����;`�����*���.n��ˋ=<yzJȎ{�7(�����E��Q������</�����K�ʍ��<8mm�������N @yN��z�ɣ�p�۷�oR,C݌��97�&��$�L\�m�|Q�UǤ�+��j��09XlxVHYEB    fa00    1b30l9��-M�t$7l�x��]�ita��<0Y�Z�_�D�G��L��8F����{���I�I�V~jZ8uKj�Lx�ZA5���Q;�Y�a�t�L{j֏� MEy����tNp�)��1��¹�o�i7(?� Q5c!*,���"��h-��]�v�Y;`�Dc��48��j�t�x�:$Q�i�j/S���h��\h�����a�ۄ�m~��R��#�o��'�u�0���~e�YT����AA6�P��� �ӵU�NfO�ɾU�� #qI�Y\$J �1t�96��WKSg`��J�:A�-_Ij6c�px:}F�V��5��Y��0]�J?\.ߍU�c��S��Oe��f1d	��{<A�2�N�r�z su=���=��#��~!#r_�|�q8�p�ˡk8H�a]�4y��\ۊ���B��L����sb��Y��r6�	���I�\k(t�߈?�p��yr�;������$���o.|����fN\'(J�ejI�x��/��Q���y�U,�,F >�ҁ���d��U^���
�G�&A�q�8��{�T�4<h^�>}o�=З@8�����鑒pm{����!"���B�T� �~g���=�p��s��qq��M�����B:'z���G�i�C�S�v��k��!�}�m�IZ�S��ǈF9h� b�}�}��w1ߢ"CP<�����JP����ό���z�V1䈢� �:��$y��@y���L�i��+1Q�<{�{�W&��XV��%�V��{�PB�0�l������]�������H��a���Kg��yk��1�ٜ�,kw�Bl�`<�;m���~ͱѵ��Sg��5sPN%&��,+��k��11�/J��n�q�QRY����(p�
�錜<̝mv�Iԥ�0�߫���KƬ{gy޿٠ɲ�pl&0��y�9�kt}ѐ2��ו�T��s�[�b��Ԙ
�~��)�&{6*�r��s�}���>�@�����\��bd��c~?��^� ������p�4
f.�J��v����2��:�xV�&۞9��?��t�P�W����I���D�
\C��.��!;`�#��o���$2�&�)����,,��Q0�C{�۝���¾T���N.��f��0�]��F�WE�4�]�T7�tq�~��`AK�wյL�m����g����3�}�7Xm�D�������������� �w!N�`h��[7+�����\Ѷ��Si��J��.�ڋ:'cQ���X<,�ڒ��a����B��s4]KW��:�fF�]���&���0&���3�b��+�����i`o(�> ��*#�Wx���X[�&8.$ɟ��]���xh)��Ъ�!��!�H�+��i��n��!������7%��A<L�Y��S\�ǣ�{U�Y��ͦ9| 
&����hx��~G�J���|�#�J����;t�R`雟Q�	����'�Z��Ȥ�Z&��)����J%�c�@T4�8o�G��?+�;D�Vn�l�Tj��x/ĩb�+����H*W0'��6~
T8=�l�gGEF����1H��}��'I���ckc;N�A��z�#���L�(�x:E�=P]:\(�jT`˂��!Lt~Yx���Y�P�<��&�ig����F�W�.��}yN�:�hd�ѠHi���0�Zfd8�uSu�R���S^���nr-<��:�����ӵ���/�ܽ��z"5|b�'%����zn���+L�=�6X8G(|�a�
�.3E��0�Y��b�\Sw�>�������lo�������o$��������7��¤ 10*��a�^6��
�m+�tY�.�"� ��mˑt��c �p%�S
:�q<î�ZP�y"/U��a�l�#��D��=R�A�B�U��h��N埽T�S���p�luQ�E�4������Y���Ӽ�/�i�r'�B[.9�	��j�O�T�S��6<�\v��ظ����ö����k@�B3���=X�q��P2�HUzt���2c�S
�����):��{�,_�K̜��4���N%JI[�����j3��ol���>��A�[!<�.k��4ú8AJ����[r���şȱ;w�l� ]�|����\�Z|�#w���ɂ>�s7��;�	ENǧ��5���[(8 j|�v{-B�"� Y�`$A�<r�j^϶_�;J�d���ԎY]+B2q�Fh�Q�?��7^���u�#���i��n�1�<*�ׄ��ͬ;'��;J��\����<�bSo5��/(  �)�Af{,�����L[O�^�g\�1��h�9	�ʵ�i���`l{�����iN��u�*qY�=�y���~���oӮ���n)��@h��[�oQl�Q��*��\�A��	4� k��%Ǡ�XMf֟ӟW�W�8�8V�z������9�ү9���24��҇�}�!״jI��˅i�O��o\\j�����ط1.0�mQ:V��m�e}��E
�����6��X���I�����4�Q��vZyMz�1�i]��iA��s#9�Z=>���I��h3�3r���0����!�4E-�\�4&�VN�lP�'��"�I`�\�x�!�Nwn���M ��ܤ��[���1�utz�y��F��Y�]O׆|���xH��_N�^>+i7X�s���\ʑ�<�&Eq� ���!���O���DUb�ZaU�%�m.9�Ⱦ�mk���l�C��c�P�e��͆ kJ��7�S����]�,6�b�1U%�H�b���-��$���u'���"�k�R)o8�`��Q@��p�{�%��Eߋ|��Ur.Cf�$��Nܥ6�,�����.s��"�ߢ���R���	�HS��@�7\p���%>�(A��Y��X�O�>�Il����:����_{��Dӏ��F���A�_5H���>Wby��dh�|�����|:��S`x�^Rz����!j� �u��!.����vI��Q� -�N	�-bY�j��ޒn��?������̗�G_�\9-���=ǩ_��đ�;ԉ�c�V����On��P9tpq��1��6DM;�
j}F��l�x�I3�V�����^m t?�$��4��0�{: ~�k?��ΐ���EbpU�qqvz���T^�쉕򼏗�z@Dsd�K�=�f����f�ƈ�=3SX����a����CT�܆Q1^,��:6�Ȟ@q���A���Q�f�t�$9�����F�˧c��6X��Y��r�ߟ�|V(�Byu<ѯ�����$�T�~ҡ�;�ս"�1����W��]b�t�`��~ԣ A�,���� X�3g����@P�$�;:�V �X�І!=���Im����&y>L�C0��b4>��qv�ٹ4[S�	�c��=�@c�'�2�%~�'�X�.�{�麖�O�.c���c�뙄-�ɝ�\�[�O�W0�U�Lѝ$ B*�}��� ~|Q�`\ǌ:��ޣ�J�68&���GnB�]桂�摧cBc�W`� ";��جmX{Y�`�l}%-����qZ@���G���".T`&�ߔ"i�o��ge�7ʓ�R��6\q�Y� Fu��6��5���\��/u��p��?f��&4�X������&��Z���V�38��y��|)�1���dVx���}��}�?*4�S] �Q����2�`�Hn���G�t:�w��|^v�y�R��eX�u3�������_��+O��:�� ��{TΨ9��f>
�ڕ]�p��j��K�q��X�Uؚ����=}�:���}xxg
Y��LHR�ú���<�4��N;����96�L=��z��l^�G�N�o|O���N~���:�$M�[M�l2{�^JT/3
�a::*�Txm&t�:�o���m&��#�Qg���U���ˮ����U|�MoI\Fb �P�	K�0�j��hUqE���12�����m�;� 9젤���-4Yq��e��;��T0�:�D��\j��r��M�m����������;�G3�b��9���z���.z�yQ?Cs���[ULu37�Ɓ�@,���)6�|�5��1Z:����:�������yt0�⵹+�̔�'���ԟ8ӜDn�2b jDT�g�9���N>p�H��5!�i�5��Yp��g�ʢ�znBzJ��b���j���i�ݪ�}����:�<'���{"�:Q�
@�5����Q��5�&���� _��R����A���y��`u��x+��+e3��DE������'>y�d'���zia��� ^������=&S��I�E_x�u��J�p"���#� �� ��j}�<�0��Jd<a�&Cgѫ�sa�wH#\1�=G7��*�Rq�+
��3F�oP���e�Y3~���s<�a���FQH�U�7�G|c��ז�c�^[�u���W�ϵ]m�������8mkax�.�ŋ-���by��,�o�Ӷ@;��-�i�V$��������x�9�G���3�9~v1�9P %$�o�x�}��d��C6`��-b��S�b������2��L�3�~�ηޟt�6"rp��ț���N9/��$��RF���������n�4��\��Mk��	�f��M�s�f�Ŝ�^dP��eGQ���n�Y:�3�������x�_d9I�\]��V���uݸ٭�0�N�0%�#Ȧ�%�>o��]�;MO��.��\��Pv��I|��&FdH�m?��\s�����g��`�Y����ۨ�LW�7�S%�/_Q>�/:��5o�����ߙvE�/x�;6ܵ^Q̀��5�[�����q��A@�Ɣ5��y6�ú6��#�B�A�Q&ƍ�`#�B���%1L�a��v`���(�ۃ^��=�s��
�ˮ������C��\�\�=x4�!��Վ��<��D��)8e����x'��R}�f�K��X��c$�pc�W����ݼ�r��G��p��`WR�։�!�}�jrB�w�����,�0:��*(~aQ�	I͙�,����
R���!���J[���J�x
�XL��d��8�믂�S|W��O�Y(���r���gNH�������\��u ���F�W	�*B�Y��$^�I�v6���h�B��v�FQ���ҹ-�T�dA_rF���
:����xO#a�>��d�8� ���k�>Ǣ%;%k{H��?s�7��=9�	0xO[�_��',>���ۭ�Y��?f+Ҧ�
	4�ΈF��l�irv��7��Z���ׅ8Yg$�e��&-c�q�zv��;�:�XVG������[��v�"g/�1��E-˾y4XÔЌ��tR����2	�K�l���!�q���~����Ȗ7B�S6�O�g0(�6<v��`E,J��q�|HO��3QwQ;O��]��Ŧ.ѓ�uդ���T����HN1?T�={ܶa�d��fӨ ZX�t����MT�f6�#	�'3g��ڍZ5�U�h�dC���p9C˷����)��~�驙��C����pAv�1�K��T%aq��V}�|=��L���ŰX���b��4�R ��2[.��T׷�
{8Os�}<c���γJ����o;� p`�'X��`����h�AM]�[��U���'�i�p������C���sG�(�A��K�'��˰#o���k�0�#�5�x��i��q�����N�ɴ�k[���\�1Ǫ{؃������#�b���J��ٮ,�BҤ��-W��ۚBʬ��ݷ�{���!�*	�۪.�u?sC�����DL9ݯ:�<�-�[�)�z�ͮ_����wH����Y�om�*�h����)\�4Q: �7�ǲY�Ƅ ����q��Y��w𼃢�_���T�>w����ǽꡇxs۳���=��	���{��ƚߘ�4N��&�����~O2��q�l�� �a�٤��V�ȧ-�i�4�>4�A;Tu-��eL�Nn���K�=f�s��)��X">�a����2܈6r윻���oϫ��x����>��^_C�Q!�Rvs�@�S,Q�#&,�2���j�J�K��y�F�;P��sPSiE���>F�B؛� Ǽ~�Ś�M�R�|ypx��C29�L�^���!1�j��/�7,�8VYM�ۂ)2Ir R8��%;�.�!ߪA�U
�/-�L�� Z(�"��;�b>'�?�4ۡ���en���ݷF��e��\�M�4*DL%)�ޜ�j;^����������ez�9�\E��5/�G�ɧS��2jڈ�8����%w4D���!1�e���Q�^`Ć������6P�MgD`y��p�z��4϶�	�2P��ɀU{-0dI�G��+`��֯�f��x*At��-[��n�૛���Ig�� �yt�;��A�O�rϣ�|��-q�#t��d�H�K�c:�(�{��A�PP{}��`��i_3\Q��v!����*�z�'t{����W����i��=�Z�!L��f ����m\8�k����IVX�#�ʆ��	�Ʀs��EIqv�	p�������aWˬ�Y`��\�	*�MD8�����l����C}�o�5#%\�k_k���m�r�9s��_ȧiu�eeAy֫J�MU����~��!�����)t;��5k[���� �߀	��w��S�n��D��<���+�쿋���? � ��:��'s)�VR��1�cc�!v�p�s(B�T"[��f!�"�"�྾ذ	�3�`$�ʃ��BG��M��i:S�*ᱎ�T��5�"�V<�������M]�� m����S�t�	݀��TK&��Ғ�lc����{��H���G�5-���)l:˔��u��#�3��s�W�º`�@q�oM����-�t��a�R��`�N��%U\�r��l��t>w"�:EۄXlxVHYEB    fa00    1950�okt.K���M��$�/�Z�vu��jPu*�%��X��tǦ$Y �Kś3\�w�&L��O��II�@��y�8a�[-�r�$M�:����j��������G$҃��J)$+�+���sQu��
Uc��f��:�0�L��h����r����,��
��Z��i�zd��5B�:8�l	Ő,���+������Y7������$��TY3r����H_Գv-��g��N��6����Y��/�Y���k�PkƝ�i�b�]��t�SfodV�=�iRT�UZ�JIV�=O���n��%� �i&*��Q C���ة��\P��� �hx����RYj�4�6����a����]P�k�ο��7X�i�a��[-���;�h�1c�5����*Bi�H�1BuwC��c�&w���Y+4=�U^��`,��X%^����^�Z�*2Vz�5���ۇm�zB��8c�m�����;D�I�Pa&�4R���bӪ_V̤Ss5'���,�����Z[#l�ۑ��'^�Iu;��[�Jix!��^K�C^��%S��9J��ש�4��(e�)J⽪��̷�Y"9Fm�X��Ey���T�r�~�4���Mݯ�᬴V���,��dߎ��< �ē9	�&�Sh��GA��\߉&�Dpa��@�mKǒr؜�N�W��)���웰
��I��$F�ҋ3��"����ei�Qpyb�e�]!1)U�<A�m[��HbBG�|e�UN
CuE"�r�9	��'���ĕ
 Y �\5��I�T��b|>��~%ǝ��.�+x��FL�#\[w�� �+��h)G�G)��SH�ds�� bm�Ґ�b)�Y�\kN�E�Ė��L�PP�-�+k8��u�
ln� �oH�hR'#D).�����a�^������,%~!2$���c:݂,����H�ۅJ:��˱C4��w�o8��Q=�_;�f��#	V��_1�ҿ�P6%�����jM��}.������t�!EϪ����ν�j3���-��c��1�6����Z�JJ�S�J�q^RG���dw���s�{���u��6U󐧝_n�Ώ�5p;���&�S�n����0L*3`Z�yf��>kܢ s��\\����e,���_z�����.t���m4Q:����������ts�:������mcV!�#�l&�H-
�p{ߣP��/mNu��Ѷ�ak�2����J�P��CK-O8l�/�{\���j�w�����)���_�i�;�M�Aq@P%(��ڕcZ����9�����pJa�r���0�+|�8 �ݰ�="�A(7��}�շ��0�Z%�r��O���g���2�/Y(���Ƽ9�b�W~J�AэSq��0��U�}��F �B��u��}H��]�)M�cD�;���8P#�x���Yep�w`�	�*(O�R�_����d ��Љ�
�!���U23�����Verur�K���lO6`;�h�E-��vб��J[j�	�$M8�i�T+�
s�����ٻ
�%��T�Mŭ&��'V���cs��k|�N��\���?������S���caSuw��	�.�CU=�W��tRZ����mO ��Y)"���Os�؅�%�61=�;#p�
�h�0ӕ+��4����Z����z�<��/ax�l�0X�nu{��>0x?�����p3��j�vu��P��ը5��2�Q�d'�����'B�����J��o0�f#W�w� �&D7�"֨�l�Z�B�ԭ؉*��v'UP)~���?A���E�hkj�K���8+�F���i0O�C:�nXVTa�[�+���P�m�T�<Q��Yo�a\a��x_P��ςW������w��(��Qs:g�� @�J+�\���7m����Ɉ��z�:���0��TRn%����1�������v]w2�G,�1H�c�Y�O�4��A���{v�����R���mC2���UOO����`�\Hޏl�zYy�wl6ɉ��d�x��qʢ;ѷ8��_ Ј'St�G�o����-syb�<q���@v\v�x��Nvy-l���'���mz���������I�tv�Xd2b�A�ۿ�G���r7��G��OGj�"@Y����C���w
h���N�E�!�PTn��g1��w� �R�� ���_(Z3���YBi�x�.��)����)eV�ر���֖��gzTh�h~�A�k@�c��kDQN�\"���&~E��w�����ެv��W�V�~�o>���_���)���&���<k���B�\�j�EA�cL�l�N�1�|5��a_�|��.C*�%�a�y֬�M�r�F���
;# ���ccB:m�
2p'^�HS�вo�SA(�2YH`�P��5�z*��1��0�<h��!z�t�ih$���~���B�P �����T�.�O\������	�)���A(l��A�- ��l��^;향�z���8�Pǖ0�
�j(ܶ��S�9�Y�<)VP�}��螅Ϝ\i��Q�a���
����a���_?~v�٫-L�����sH����){�v}=,K��-�~���tc�,M���i�6l%3��2�(�����Q�͠�1($��Ҹ�%��d�k��3
���&Zk�vr���y���~1̀c%��&5 �03����}n��F�3����Ă�Y��M�;7����RH�������^���p@u1;�n��x@��t_.��V���͍�}�}�x`
iB�(���]Q_��^����"p���s;tP����YP��m��1T��PS��`w��<�T���9�y�2}W@���%�ݾ�z����lS�>/]I�)d����'�2�iGݮ<����Y��U��^�������ù�W��@�=�dE��u2�����Dۢ��Vc��B:����Y�t�:[8ܔ\��K��;�w��i�įP���I�jr�s��ꮾ��ơD�{����jO�j�X�̭I%Fn7�á�bB�N�L�;��"�x�W�.nK��v�ަ�ڡ@�'� �*�1��M{�O�x�6L����v���7��Uhy^�d�O��I(NO��{�EC: 6f.�S�m����_P��n���e���~�&�����6-�J�Q| �:sh?r��_�X�����'���Ԟ��������< ��+H�@�E��l�r���φ���Q�O��B/�|b�)b(��bV���� 0~_xN�0����hg�L˕�FZ�&\? �'{��3�-E�6����;7X����nn�ͫܚ�r��r�)u�PnI�g�Z����.zW�<k�+Z$���cb�5;��{H;��3�*Á�mH1$���z˖�h�6�����syLl��Za������"��fE�[��ED�����Y�c?����0IjX"Ǯ+�7��ʐ�Y��*E_o(H�5I�A�<��ھQ8	f�M�K�u��<��� ��x�OOՔ���W����̱�_2�ct�IƖL0*IB�q����M0�#�x|(O,�H%нi�\�=и����5�@�R'��%�I\M`��e�s}?R��ޜm�qkh�y�S!��w��Cs��9��~=Mz�H� ��"]H�4����'�B�2�mt�a�wl�햖O���TW:Ŭ0	Oq鿙�}!�T�JS�eN)��k�Qi�qU��B����0h,W[f�?�*~���ط��򔿉�P��;E�һ��ˣ��>�nq>�ِ�F��d�4-��wq39ލ4�GLg����pnz��`�ܒ�`�~/d&��s�~N�������e#$����^��C<���=ێ�V�pp�ko�-cp~q��\T6��4Z���*�9.��IŇ�9���xJ����n9����V�Ѐ���A� ��4j6�O'w4M]��S���<\��Hh##�j���(���.g��l!�JR��1��� �|�z��ti�V��&�� rT��=8�ѻ�e��L]��'��D[j���g
�S�I���Z�L�p;�}yh�~�B�=��ڶm�\o��ڰJ�*_��?�WoYBe4��T�G'�L�'g-u]p!6��T��5zs{p-��-�����J��8`��#�'?,��)$�Vn]��f�
"��l��xB�F�<|I�=vf�Ksƍ���=��Ea#f!|%�� h ���K�<�7����q���Ú2p�*���km0 �Ku��jG�_����8'1f�L��^*°zݣ2�x���`7o�@&�'���b�ަ"���K��V��(?���G��f����y��$�p�c�����`��El�v:�������cfrK`�!�^6S����f��2�Q�*I�Ed��7�/�+П��bq�g�$���+VQ���z���Dpm��AF�+a�#!�����I^�0�e	^hG���c��due�{��?���/������V	��t��Ni��1�o��l��I!���>?58�2�����q�Wa7�U$L�c#��^;�5��YeL̬(U��-����S�d�B���U��	�u�3T?�~y7r�%��^AW����t� ��5J���>@L1:S�Ӂ�f��[4&I���i���sE���xd����m�b���'�M�#*ӑ;��ﬅ_T�Ul�%��ԫ�I(3Lh�����ұI����#�4��
�l;�h�#z�Urޚ҂n���9^����u�d��9A�и�q�>�9&��U�Cy]
n�z�w4�s ��iw�9V��[K�~)�Ep怂u?1T��"�?fŬ�z��iw�w�|��a��/��nL�W\�7�ma����-�����!�\�uL=�l��u�}�+|m9rFʑ���G 0�^�)�h�|�~ۚ�t�ҥ�K&�	��E��\H# [fP����ccM��/a{���MUx�<�@\�@뜟H��]R�$�-�ƥ��K��������MZ���Ȟ�]V�[jLMk9}Ep*�h�tn�V�H�f
��4��w�"b�T��k�·�]�0�mh����yKs!(���뫠~���[x�\�:�3=:�P����5j@��mr:��ު���s+9Ht헯��;p��e��hw�x�|�����B�	��{�E��g/�8���B�p����P�*2Z-*{�/^T!<��!a���ký=m:	��<�c��=l���\߭�҆i��͇�����Z���QX�Jo�({��Mk��!:� ��Rh{�7ݼ �nDjC���>��؎�����WE��:�lD3�!�8a���ޏ��M����s�ǥB�� ���`ϰ�^���e�B�����W��$(ۄ���%�� `��b�˥FTG[|8]B\������h@Uѥ�%����<
*:�ֶ��]d
\ȸ?&1J̌�,�I�(|#�GH(�_#5޸��DVs�&�f�SQR��2Ӿ���ev�;5R
�E�D�_P��`�W�����ܮ�V'�7I�<��)��YC�9n0۸R�8�����Q(V�U&P�t���N�I�qSq�(�	�}<��)�5N^� ����򪀝A��J3� ��iQ!�m;�IA�l������8^F`r��
��-jYR�����w�7��\�ς۹�}�gU�z�+Z1ݢ�&[�/�$���Ύ�M����>�����!��et�n:�܅����l�=\aڪ��h��-'�k	���Ô�׎c��~��4�q��3�D���b���N(�#�H��d�Pxb��]Fɣ�OmZ��C%�k��]D�a�;-�9G�5�����̩�l�p�����Tk_mT���$��oV�^_-�ܳ����T�/�:n���Sp��,�j��Ԁ܏�X+�w�v&��R�,�קV����;����pG(k+!�r����]�喝i�X�W����q�=�_/\�fX2R���^���_���h��2!W��q9�+�>*%�S��ʧ+�JYgI'L��	0�g�3Ew�@]���+�ɨ�;�9�W��0�;u�Nm����:Ԝ��C�6yL�+�;K�{��$nvu}��[]��M�;e f�yjb|�����Qxd]�S���F%�ߍ7%E��9|��c�S����Xd�O~�ny��R��u���Z_�����P�_��F��E���eS 1��i��M���W�1��}�|:�N�E����%P\O1^��7�4Gܫ+�͑�H5�A�?P���a��n��g+�D�N��r�~�F�_�M�`��h�%��B�aR�V�G��޹׶� [�4��7�r�Bx���v(��C��
�ϕM���eњd]nkǤ�Hs=M)Ы�w�2���:c� �~��՞2��C�-�-E{m5uJb4%9eIΟl����k�Jr<�v��,�ī�X�XlxVHYEB    4f27     d40��`�E�,y�}Ǵ��1�f
"�LQ3X�dh/U�x���cXۺfC���iA�e^��:v��A�d������Ar5)pIX6nQ�����B7�����
�.�4F��#��f������11GM�7�=/���Oߴ�K�����qs��[��&m�e%HZ�煘QO�T�c�D�iu�,���$)+%��I��#�D��vO�aQ�� )70�F�%?i�2�B�������V�v�����A�T2�ҴH'�9B^���헛����-�T0L����``'�#�6B���9K����)�v��l�Q7,�Ub���z�,�8����~�N�Y����Ǉ�0��~����x�w�R" ���x�i��0�m�!5✶��6������0S���0�ٻjA@�ʒ���t��sp���
ψT�-����;n�_3��'��[�U��{� ���'�E�s��X!��-�*p=9tSe�E����zV�3<^��h�����)����K��tA��:��#򳵇�d�s���D!��][���'��U��C���[�54���惜�I��o�U�:�;ɧ�N��f�KmQ	����r1�K��P���=�'W|��H/b7��w:����M�\i킁��q��:j�V��Y�&�]_S��d*f����nvx�3z�*aK�^h�/8�G��tt{21�����p!���Ř��!�#�����KR-)�U��*6�̒&���0��@ٳL���Eb��T���/mZ�C��wtTy����
x�s�.ˣ�-�[(�:DkZQt���I���Dk�B�^Ҷ�Oé�D<���hQ$B]vZ��t��P]�ڜT���II�Kȥ�Cׁ���Ƶ�8�aQ������$y\����,�kg�Ɨwє����s�@�"��"'5������z����oT</+���Ņ�03EM���|:�h���:�1���O�,¾G^�O�����!�k�+4,�S|}�Lܘ[�)��Lt�+���8�<�s���BGd�.Q����a�9!Cw!������K�r�~h
�җ�f����DC�5�_,38�+5Д�2���R����R��x T�e����#�����$�ߡm�������k����r���i�� ���i��� )?HX��ǽ�5��eR9�X�_��I�����4�4�$�S��?+�ߵ:�1⮝��
P|�����*�Kƍ�{��k�vV��M��P��}������������C#�znf^���#�d���㔑fJ��/ٰEd�`ȭ�W~�Ė�8 ��'%�&����_!5��4Oe;ʎ5��*d�>V�$a��h�#J�	���"g7��w�E��جJ�#��i|��V�H�~\����
=���~�s@�!�/nz#H\��܀��\���
̜#�fxv��<o=�E����ZR�Ȓ~�R�AT	����n�)��|�xI�Ή���-�\X'��x�);�C����0�����F�+��#������C�Ȑp^9�`�4��X�$��)�y�I�UI�P�ߤYoqPjVZ8mz��������Psz  ��+������8煾���{� ڌ��d�rQ'xN�ݧҥ�C�a�z��ز{u5����5�c��)܎Kh
I,��&��R>�ƫY?���w�%�p�2'L��xHǑJ�zD�+� �	N�T�Y(������`�� �3UC�X����Jǡj�ڞ�r�)ߝd��9�pxbs��������պ\G�8߃BR�H�K� A�������m���U�N�
��_�d�R,?�汄 ����m��'T�v���}}�\�����k��V�ze�{�J�WW��tJ=��m���6�)�o�1Y������d�>;������h����y�ʠ�^�e�᥷p��O1|��C7�@��jMg,��0
Z7�jt7�|�.��˨���=z���	���'�:Lя",���aF:~!�=Pm��բ�)����n�!M^��O�����R3�X�m�09��b��r��8J����6�]`�f��4ڐ�-#x�dϴ;�^�#g�!��"~W���`YS7Ξ́��	�_a�� bH�=ls�\@��D1��b�7�G���o����_�Z�[bJ�>]����Ne;�	�J%y\+�T��CRY��㹛�v\��"����MN���� �J��.0�- {}�?}��r	jd�"[�T���z��.�hOc	���NY]-�-��f>������o<�<�]��vp��UB98E��'�j�rOXt�u�*�J��`��D��W�9WUJLL\1���3��:��Z,�3jI�ک�@��n�D����/�lJ���®ng��k�۷�)f����#@D�-�v��-´��h�5&1���@`�t�@βH�ܪ�!I/��7L8O�$>�'���Nm�}���4cF=���H�\��<��,)����0�}�J���EAM�w*��~B��5ʴ�)x~SS n��0)�!���T��Kg��?��5�f%!{��|ލJ"�Q�<V�Wes+q�l�cА����l�\P��������/��5n?�u�N%�IM����+�E�6/��fE�SS׻���p] i�PɍF��{�I�R�Ƒ�&~;]?Y��N��8�0n�!�KYY �O�WqB����O��^i��\kE���@D-��ἧ���:%�?౹�-=c�z�sN����<���I�E�W'|=�`�K
[e��`SsK]&�{ٖ��c�y�W_M�׌'r�
��j����<Y�lU��~/�H�v�-���/uG��H�Hf�~�0�Η�P�Y��YƱԻ���]�PFD���F��t-	���
X1��}�C�0UgWM6�Ve��E�͜&r��v�=�Pe�ZT����Zy�۳���-�|Ҏ�E*m����}�CL9*~���#"�p=ܙ\rJGΗ6	zn��ɭ[{8(�����4*�h���ww���`�S0!f�{`b��j0����6�2d�+����P�NuTÇ?EV���Y�y�'���I�!��Wa�椀O$��<�,�e�j��9��P?�>Ͳ�UL;f6�M����9ˏ��eig_�H]�Ґ܊�}H��O:���=��������l��n�����m���̒0H�+��0��Li��*��s|è�bVff&4y�2L��������ف"��l����ʾvx��Pl�b~�w���Sw��<�7yy�?��ޕR-{��&m⬍��d��\��I����f&^� �� ݀��,bf�gvҏ�����H��;�[u���x�+z����X��k��3$��2��(