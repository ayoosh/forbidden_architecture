XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ER��L̳aA���� ���0�q�&�H0�����O���+�+�Cn��Ҥ��dz���햝zPw�[���|�� u�ߐs�rDfTZ;b|��U�8����zf�7�\~[ݤ*Q����zZ[��H��IO%x���TKŭ���ʠ`��6ʍ����|�ŋ%o^�Qj.L��r����S�3��\O6�x&TX�������{�	�R�0���
H�x�T/�(��e�_����1]~Myy?^�OW�h/��4�s�T��I�>|7�>��V���U_��re�l��=\}7e{ҹ��ŉ\ƨЌ�"�>�N�1������I,�����g~�m���U��Q&�i�k��5�TP�L\���(�q�����Hzr"��v	�Ȕ��|��e0!7."o(� �����^����0ß6�cכ�SIjL�wVx(����:�Þ���T�����#����L58�7�B@�X��[�+�R3}����c���	F�}�Ī-]�H��aā�d@¸q�ѝ�\([k���~���Dlhi�/@����	�f���-A��ܟm�t͙���,�-3W����?���G���=����q�S���LD殮bȮ�@k���W�ËiǓ�����j��ji�u�׸�_n�&�}}+���u���֑�z'F~%�5�:��p�t���4�-�#�a2��ݣ�A.�n��_��^]
<��vo������1��E
�V�?�����ʂ'�K|S��6���4��0�L;ԴXlxVHYEB    fa00    2d70jvbw�=�)���f�?	_\oY�6uu�Y�*�p'�b����_�A[\3��`�
��6�zԍ|4�_�aXҺ ��&x���-:C'��y���e���Z0��ar���%�R�&�Q+���R�U���ߴ��[f"i�oXhK3�-���I MW����^��	��>�w-���H��p�5�T@G��Eڞ�3��ȫU������=�b�kQ�|��p�Q~�x
"���#���<c~���`{o��-��c�����J%v�w��Ӹ�~\�
?��7�D1���y,�dlO���Z�W��*5�F����ơ�u�]NI��}��㔐q@_�JLS�DӞ���Ѻ��k�	J��H>����1�5��2�Q}P�������������]�L��4`���s�< _GBU��G��Jg���F�h�?����?4�t��ůSaZI����
���k�]Ɩ��x�+=�Qn�U0��E��Ĥ3Bb%�ؽ�0� �04V�>�8�P�ò�:.�F��΍��g�$#$ZW���K�e�B�N�^X���66�5�(�"�f�x��k��50�?i}�QCr�����4`}�BE�Ɗ`�\�"x���n/�B��0��bt4S[�4�I*���C�����(� �����q'�k�6�>��JWg�mS �g#ј�",~�����۾,�N�J����\SB�����}�$=���]R�C��a�"�-w)t�� �v}��(��^��Z�G"^�+��-��g|)�e�nQ�K0y��˞����O>�B��8�x�	�HC8WV�G�b!�s�g�9f�#�6��M�Iq����r����h�u�~9�AӃy�:D�iL#7�Y���+e�w�؀��xޕ���������43��e�K�b��|@���dM*�p�@Tc:1��	I���L�n\���������~�,���ݯ�f�=�7M����l�b���p-������}<Z�̢؎��h?{��*E
E�����y�m�ǈ[�\�9����3�ǖ`%sv�e���%���'��@D|�e�TY��S�[�d�EK񽨩�S(8ω�,�V�b��`�&)x=/ Y�?�+���b�����2g�}mlmҾLtu�={�!�U�����{�sQ�1t�ٝ�;�K��>bm�7�7�8'W� kaL>ZP��Ǡ��\(���RR\H���-����Ɉ�9�(��l+����-�ڧ)
ބ8GfpG�Υ��AӐ)W��n{F�)�lǛ�9O�r�7��$�Z%������W�VQ�c��A{X,\'G�A`�˴O|rRe9��t�\�G���^G�Ǜ-)�J*�Y��xw�o5��䵦r~P�YZO$�L��h�S�7���>�H��4ᑠ�*~�9f�	��$������9mI��'�U{?��C'�f�_Kj��eX�u]��=Ѫp��$���v��&�K;��"x���j�%v /�QN��y'��n#T�|a>�����>O��'!�H�Vͦ	I,7��ȗ{����̧ٖLFQN�J+�Eh�!%E��Z̯���#q�� �����s���L+H*�	0�Ci ��{��\,��X�+�b�{�厫<�h��6��U��y@��e�CWQFaKG���h��~�!�X!��;*T3�ɧ��(E����̳��v�^JfF9��LΈ�=F�~�M�7@�ϟQ���4��B���<�	��<ҊR"�㴻������,�oC�K�˶\���C�L��kg؝D[�1��F�e��3Kpf�-���E��U�]��:���_ӷdХ�M;RZom?u��WH�^u�O�,��!�͛CS�~w7O�t``��Y~U92e��*hʕ�+�;��UΡװ��C��ʦp⹻�-�1|�EJ�zR-���Qg��l~��|L9O�����s��t�C:�/P���5��x2�j�A�u�Z��14�z�k��� �D�/B�1���J�p���gM�>%6��Ha����.�+���J����S4\s��L�L������:r���L�-g�M���6��wh^�+D�yx_M(#^
�����L�џ?1�M�i���B'�)��Ԩ1U��0;&����x���CW�b艩x6�����@OMnNh_�7J	M7vB��e��ufB��:�[j�8�خ6�w�J���n'&cN����e��l�d/�cϓ#�{��y�e�$�z��٩�	X�|F�|�C���GK�<�r�:��W�/�������Y���3H�H�]y	KM�ޞ�d�^�R�=�|oQBIE0%z@ӒX�AI*���'��\T#y��?��&Ip�m��/v���'Y����mh�����MO�nm+��"�Mګ@Y��q�4��9�AY���z����$l�۝]4
%}�Y�W���rh�s,p?.3G������xE���9��,�eaw�����"��1��/W�L���o��t�1�ȅ[�
��J�������c���Q�-��4:!|�8�7�wO��Um�ШMв˘@rR�����n܃"����(��I����l@3Aneti~����Q��(1���m���uؚ�-�i$���Җ+���^ԧ��s�}uB��1�`a\�6������_f~ܐ��a�|��,h$���(�6����p |�l�NQ](��wx�B}��S��5Μ*�����L�b��}�1���LX9���= ӽ}f3)��(s*��f�����,%Sв�j
�JeUG�/�CC�x�p}��N�4����8�2k������o�*P�DK�(,�6 ^���m_��J�tț�r:f������pD)!�6��{<y���{�I�#0I�(y���5Fk���^ZF�>>��_�Tkז��{���g�E�w�d��Z,x����uk�;�E�'b3������=F��[l��އo��t>�G�֕�uپZ3'p��vî�u�n�4t�bё�y�BG�Q�bfan�~����i�'��9�C�\�P�G{s@:[~r�wi�$��nZ��7��X/scB�J���3s�J����D�,��f��,�:>�F輍�;�
;ĝ`?�΅�W@Vv�՚(�Z��]�=��rȴʷ�%ı)>���?���%�hТ��`�� �:t�x���Q(�Ϣ�7��ҕap�[ ���c���9�H���hd/T���?�9�ϋ��I���,	�/�kc�#�E�6����4<������Dxtk�J�͜�3� ��U���4E#͝]O�`���`����M��v�,�DLE�A#�e�����&E*Xq͋�I��l͔�w��μ�b�U$�m����j%�Š9~m.G3hT7���B�=v �ćsj������~|�j( �H/��B)�`��y/�̷���\���0�U���3��T��Vh�#-ŋ$A��/�)va�&�#j���caI���U����*lv#��4Юi�Č��6U���vf��xw��T���[b&���j��xK�U
�8}A�nh�K&uo������
��c�Q!2^�Ƽ[�*��V�A�d�#�MH��=;�^�NAc4gYz	��͆���ܫ�ڊ��<�r���Ĕ�2��a@�bE��{��ܽ�]���ɏZ�@t���Xm;?U�2#H#ר�x��C��s��|�S.���؉8o�Go���z��Se�Db��ݯKCD�y����Ċǫ����{RS�.0He��	�!NU�4S�Z'����okL�D��R/L��	��E�.�S�7�6���anF�F���,^�,s�
��o*�J=<�,���n�	�äq��\v��9�緯kAc��%y	���_e4
}��Ii�c�Vk/�S�W3\�ӁK�B���»]o�����mJ1��ӻ�4BY���-(������',�P�*���e��HL�W)z��P\B����O��g�����AF��IX�Ҳ�}��4��<��H���'gm6|TX^�1Wgv���S��H�JKb>[qoO����Z] ϊB5h�~�J�yb�M>#�$\^�B��KB�.PY(�C�ʒD�.�]C����Ĺ��,aI����sY+3-_ �.��H�A����Q�����91D�p�_k����iL��f#Ӊ�R������>yQ$uoL�F�&�|��JZ0[��q
�%K�)�������?፻7C����U�d$�q>;b����ε��լAv]%y��0a�A<d�b�f�??h�'�B��%Sw�5^GBD+O�i��n�Pe�Tt3CTJY[���B���4���>~�d�!<rŧy�CC����N���T�<*�BcL��h���v߁��-����uS(�C� ޥP�5�.ja��o��z���}�AC��ϵ����#������[�|�,w�ټx2'��8U�Twb��ʶ�VQz6>.9�-�_J�`.����[0/O�������n�8^xHy\ĎM��y`�
�P�Y� @�7꯿�/U��������]����M_&y6H�xvz�Ր���:,��^��6K���^囇J.��IRw��A��._�DK�3�&���WX׳|6����qX��&��Z�c���N��P���rVr�=�R�l���C�ع h�z�~Z�%�z>�o��̗H?�~�5�d9�M�\����۔�b�]s��+��*"�y 5���d��V�W��nk�D�2_�Y�v��e�a��#6�;��Dg�=������"�Q�4}�~�c>T��;h���s>X�?(�G+ ]�v��p�]�]�|X��ȏ��y�_B�'�
<�VG�ŨW8�D��rN�3&���}�2���e��8uC�2r%����sv�ĄN�Z��n,��I�.����!��/��<d���1����	եݧ�1��7���U��w���l�^ SMW_�hj�����p}�D��|�h��&�r�2�N���^kg���͠�]����J���(*��΃����戅���9�` �L>��"ɽ9��\��XP���$��X�z�fD����2�6'�K0և ��%8 $��)p���Mݷ��5-|4��9�ieV�Xܛ�.ֆ+a���W��~}�Ї,Z�]�ǟ����M2����)��6�m�������ro|y��dçfn�zwMk�՗�	v	�����
�}Ԫ�؜�l�x7��n�Ȓ�l����ź�(81�L2�V�DL�Jq�9H�@�<�Y���P`�~�����u<����u��x��^H�܄Np���G�I��F0#������~��Π�%X��t<���a�J@=�?��v+kx��qE�;_���S��M��]X���'1ӭ[�cIM͵�}͆I��[c�_gG��n�,1����O@�$^Ǟ�/Gy�\�z{_�>w����c�=G!�q�O��/Y?��a�c�yR%!i덴�מ�E���xaN���3e�ѥJ=ŋ*T�p5Px �
�Ė��`��d�Q�S��s�~Q (�ߧr��U
ߣ�/9UC�1��?e�,�
J��R�C&��Z8D�'o��lER�KF�v�������3�Z�Řߠ:-�t�dWF�	���Z:Ѽz������G�\��� %b�I)�9�լf�"0k�s���Cڰm�;�f�?J�)�F����*ḙ=���@#�9�����xXm
�Q������J�����=��މ~�N����*�es�w"$�����ӯ�.�EP�C������S� �&��{��N3d�{j�k�]���|�m����ٻ���2Ԛwg-����n�з��SZ�����yg��L�=��9��0�n��n��	�6=A�������'l��˵�����E����K��x@����r�,�y��������]�i^ws��L����ϗ|��*��͟�1�Q�]]g��~YDZ��:�n�M��2)L��-*�`~M�b�9�}�ۈ�����l�va� O�A�¦~_f��R�&�)bXG�>�5����6L����kB��c���;;�U��C��ym�ͭ˖���n"}R�$�Z����:�0:���2:h>2O�h�T�pTm�'�\+PJ�Kڻũ�~���C�̗�N�X��v�5�-�ڶq�@��õ�W1Ac��w��5о��ja~^�Y���q�JT��yFE!a�<��O�>�.Ӷ�c�*�sW4�:�8?i���^����~�}�Ť%���H 0�2��^�Ӡ��+����L��9n�_z�P�����c���r���WU�A@��x�c7����ڲaH��w{Xk[�:�_�rG��U9{���aJ�&R��p�k;��C]�$�^��!쿛᪱�m1�_g�������J��14�%�.�X�J&�(�7CV�s���e�G{K�S�n�]��c����#޸֠�����H�੍������˄uV�<�P����ià���X�.���z��24ν��W �
�I�
�R�	����}=��5ckj,:N�.|8��x
M8��Tq��T��r7��9Σi����x�� B�hn��+��W�p|j�?�K>����_l�k��yޫ�ؘ�zb�o�I���b���ąW�z/��(o��'�UaL;4$�^J߄�z����yDƖ�1�V>Z��Ť�-��ܴf���!b_Q�j�?n%�����M\T��	��:����y��|08_~{��"�
��������B�^���~�uX�/�i�7:���7���샸K}jKc�Y���r]�_'>��vkU�-=�Wh�<�w�D�����]Đ�2%��iO�j	�I	���wiU4.UM	�����<�������r�ʃjX�JW��y���J�!� �wӼό�x1l_�T|�M��yF������7vC| =��zo��������L�(Y�:�Lxj��z�K,��И�����Ss����N����Y�f�~�[zzXPK�4�(�Dh?S�=g �D�B515i
A˧��S%%�O�/e��d�É� rI=Ο�6�e���w���#�r"^7I�>�q5�Y[)}�_N ��kC���ɡ<�= ���\����W��7�\�������X�]�$��<B�pv�=TYH�4]���<��Z��Mµ8�/�$�����'��JGV��mt�z���d�q�.Hm�P���j	�;ǳ;�Z+vc�2",��j�o���bV�����Uˏ�c'�1|����5���ۑ��C�W��n���8.4��"J'"�F����y�R��N�Xy�g�MI�M(���4y��"��;���3����ZL�h���,D�fe��7��\����t	w�5�^�x����	[�Ѝ�	~��_�훧�����܏ۄ�6a89�	0�(���U$�����~����Ld{Fҟ}:�+���
�7I[��بi�G?���~���llq�[��?�tq��yKRρ�F�z�d����"J�11�>|��+t�˫�V]�����w���~�T���:�gVά�Ǡ���j[M# _��u�o��8��@Aղ���u��0SKT�ǔ�����ﶿK�G��9���7,�4�i�jrx�;����?Jb$�+1��NT�Dp0HA�Ӹ��o����p����~��ԭż��L3�*��7����m��5z�^i19�*mP����C$��K�̼�n�w�c�/r[m̼�<#�[���M�R���8�lJw��hm~@�x��v��jR<X?��̊lVa���CZyj�v�7|��:��˂]��W�|��H�~���v6O`v8�����&EVU@7A�j��|�Sn|:LнA@��,��t����i|��8�Oz�__]�V�˥Nꓺ�&2�o�5�g��֎��������x�[�Y��H�}�o���Z�]o͇��P��Y��F�Q|�IA���S��r.�CWO�H�l���AY�Nj�T߯��)��P���02v9�Zi�2��oR�}U|/}���Qt~FG��c��1S��9"�#"𷰊�n��z�Uu�e͵e9Vd9��J�ۺ)K�58��"��y��q%�t�~�Ȩ��6��~��4l;mG�lG��Z8EĈ�����f��4�OL����z_�2�q�g4z��-Bb|�������x�2�fJް�x!����ۜ�Wz��5�����G_��X9�M�o$�4H�*��oY3�>���&�4�?��Ի�Q:��9���O�($(�ܪ��;>|N �6���р�����r2:S�HD�T��ės����٧�3#�a�����AUּ�LKj~`��f�X�wU)ë$n�]a��Q�Ƣ �	vI��>>o�w/{P�zH��g��q,�A�Aq@� �Ą��A��qB�]vl��܆ ������Ւ��ґK-��)y?'�4y�V�ߖ�:�JV3�m�?�x�Bz��2�A���׫� +�gWǰ�t'j�FV��O!��-�����.�6#������31������(.VAsI
���x������X�dpLU�2c��2j�Ut
^�7=fLR� �� 8�u�CCf~Ei+�u�'[ZD0+�DH4o�k�]�'��)욽��KX�9��L�T���V�M3$vhI_��W)�=]��&�o��o�����P��qO"g�CB��.}�]��b�[�E���!~5���q��(I�4 C�a�Fٌ��s)�-�N�����2��?U�,�c8�@{z�V�߫]!��$ �8�z(�<�kK/<�6E�a����H�h�,63@+=r���T��34֗�!@-�w>X�(-��pӗ^2F�H�4����G ��\H�(�G�j ��֍)eRXo�Sppj5�,N���]U��{��l����A3 �)'��˳��{��[c�e��G�Z1�*�5�5Q%]F�כd�w��У`&;�>��`ˎ��?�W�NC�:�C�SK�a�ǦQ
B:��y�N&�&:�.��y�a3����9�4N
�T,���� �ψ(�(hY�^�f��IU��:�Ҡ���o�rGD�<�2'˚�+k��-�/��E�%y������Z�7���ɓ	L��w�.�ͫ鿰=���z���ݿ���8B�.�n�w�ө ՛�-Ik�w0�O�hw=�E�k�s4D膲d�Z8_3��O����_W�#�����J���`&W/�:�M���m����߯��%�r��N-)%����o�e1e���;�#c/	�T�0��`,"�������.Xj�j��Є����b���JD4�#��RS������S24+�(rѸ��	�$���bI3J:=˷�Cw���w=D�����`4���iJ>��N�Ue�6i�3K�cu�'d��_�?r����7���<D�>�$�ކf��̥���UT�w람0��������T�<��k�*~ν���)E���1$������\��q}pݠ �,���_� �se�f�DZ\OP^�g'mF��}�~K�����L7��[D=�Ȯ�2�X�8���(��o�8/�A=?��;�TC_V�"G��8q�`�s�k����O�2�kԒ؎Qs�3cokxe^�x������̊�P;���O�[7��@Û~���s�P�VjI�����-��+h�X���㲥%�b��V��t�s�W�Rĭ�������8�&�8Y�9�K�2�`�3#�<��*��7�B���>YA{͔��� ��S^��~�>rf9" �!~� ���!S��]�ϊ� �����dbeP�px��bb����&�>��ZD�e)��)I�����Y����yh��ߋ'ϙ]��������}�9�;2
jvc����W���*v<y��5�ͣE�]z�3^�f6���8Z�:.��yTR4����b��@��=Ax�����3M�anv�I��U>X"�����	��H��*�����H����s�mUڻ��g����yx�B��1��L�=�����m�6�A��@�=uɘ3�B?M��3��Ё�܊�����+��ۃ�\��mL�R�\�ֵ�%`�D��f#�G#��f�8�/�^��
���fe/�M/Zֺ#@L�������L�L�0��`����ywCΝ��^��JMY�>�d�1�n�#h.�e	c� $7ܜ��� 3M�l���i1��ٛx�M�4w�;B%e�]}O	�2-��_^y�v-�z�*#(���I��Q���`6Nm�J:Z��Y!���@u���>�rX��|aX"/u���c�E�פK!E��;OƷ����l�����&�!���y?�y_��)�B&u*�Bj}I�DWz�#���MT���<�Z��z���cq~0ny�<�6�����;�`(<4��Go΃?������ƹ]�~_�E�V���$j�[V���9f��������^N�e�[�ꈠb�oc�e$�BY�dLy�;,�"A��mگ+�(gp�F����0��L&6��8�:�x����!:o&�y�],�7E�X;���߈�IΙ8u,4-������Teu�|J���H�F%���ִJ�#~��4ëѧc%�lE�D�l�G�Ee���Q�cp�}]�AlȅF�GXҎ���/�5}H����U�9��֐�$aĿ��~Ӌʽ ��md�	������R2��p�&%{+�����K����c�Tr�-�J�b�W�0�r�v�@Kt G���]�h�h9 f�!l%K�Y���/��`N?Ʀ;�;d��`�E���)v�v?}/��+�$3���^�������=X^>gi�u��BU_?ޙ��>m��Y��7�b�PR&�Em����w����H�ů�,-��F���
�/�&Ldr�$�ub�N�oߞ���g�j[*sHP���wm����R׵(W����q��s�_������bTWЉ�|�6z����٪�HgqSbLy$]�C���{�1v&�o��_�U�M��w�?�$J;��n�?E<Q�g�IO����sP��t�າ����G�|i&�@���9�E�[A�;�|�c��G=�D*�gv��[��,Xu0�.��*H�؜-��N��
9�3�a^�^<9�.g�ֶ/I��Z|�:�ڍO���jr�vCYjO�F��:Q>��CrA|�����\��D�=7̆j�P�����3\&��G��I���g{YY���I��CϚc��j�"y��2��������Ƹ�|1��` ki�ÌGw�|ݜc^  �&��4�����58���c)1M�9����wް{���^Ej
�U?�$���kQq$�ͺ�<��A Viic�(�h�r�3�z�)&��h�q��aw��GT�&�&&�Dk3(�טt��K���F�Ξ�_/���ɩ�QϞL��Gyo�ڏC�J�/��8�%f�R�}/n3<s��2wK�Z��{,����db����dxC�	�ϛ��6�W��Դ�Z���v��XlxVHYEB    5829     ef0��X�����l�ۛ���+ �C�U8������
��5�C��{��g4�y���K��%��h�E��Rh����]�]φ����K���/��8�㨤�ϲس-�A�58�*j��
��G���v�������{��N�e��T-��(�9-�7�S�N�Q�*SA��M\��㣔w����t<:��ڂL"p@B�Qn��i�<�q-oSaD	 3�:i���(��!k�`r����3Q|�K����o>f��)ޝ�9�����҅�����*t*t4�@��w��)rqi���lF��c�Cƃ�!zd5Tw�k[��ݱ���l�e�v�>�pD��%b��d���g}�Lw��!`��%�$��KE`<��#O����i��1���Cn�zkTj���#��$����W��p�3�>�oH�򺚞��@ �� �A`�SdR7
�J18-vT�;Z���"�"H�+0�t��W}iKN/��s/o�P��"��˹�ӓ��L>(�|u���
E	l�35\�����M=�&熠�	l��t/wg��ˍa� �bm��D��5�8NQ�������x�SM�x
D���$DcɚU�
����z!�4�O\zO �0q���p��_������=bx/������Y����͋=K��	�)�&{�^���7�(}�H]���@�hU��[$�؝�`Q�5���� �� Y(�40O�7�Ѓl��0�!�%�9B�Z4��v42hǩ������|z�r_�D�*�AwC��o��G�#�#p3��5*L��K8#�Ĵ�-E1��]�ilQ{�a f��_,"~�#�I����߮���*2Y*�(�Mǧ�~f�厀�?�'��ڨ[����8�K@�6x�G`c�YM�&
�l=��ڙ>p�{�Q�z!Ӣ�����䃼&��A�'�L�E�-&�s���
h�����/�|��c_ܮ����DM]w{��v��/��Z���"�_����7Z�Gf�|/�{��?�p�/%�?�I\�ɓ���!^�j��ȓ:���ԩˢ�6z7�'j�]Ԏ�K��0�^<}]��0��?vP�~�)�����U����(��;6�ՈH�obF\z;��b\W����]e٭K�d�(ks��f��?���~O��߆�&��Ҵjan'���q*�,^"}���T/w�BE�7_m��X]���D{׃lh5��h2x��y�W���%}�9L>N.��%�5�I�=A�-a0�ay,���R�6"���C	\�~���wo*k���@�q�So�($��J������ޏN�_��3��[�XH��E$<��ٮq��"Z���i��Qv9�3�1�7n&��ׅ,:B��yd��Z�'��c�6��@ՙ�Qz\�~��R�E�}��[}Wcm��HN��^�MeE`a���%˗HX��Nq]�½�ǰ�����/�2#Zת�6��H t��ھ�I_�gc*]�)D�e.Gmvԋ�¸eZ��Tvo�~�ܧ��$�����S�A�ٷqa����bN5��.��)�/H?,W+�Aт ���ڄh���[�twz�JP�M%�������OɊr��L�!R���4�H�*6h�U����)ɸ��~u ���a�Z�{�EQmLs�ɝ_c������4���� �H���� iJp��.�!/��رTP�/�.(Z{�q�Ah��ᯝ��f��w���so5�k`ͅ#���O;Ӗ�toM���2+�j#AM~�ZN�av"@�bq"��7B)�,�GG�G���)�2���g6���������v���U�E=���z����4o��b\��k��w�<y�M��G�~.�ľv��_���;w��h�D�y=�˚u���l%F`�.�&������*�d)!�q�O�t�wqI�ι�TModI	zzu�Ph.�I�]���}v}��J���-����g�p��	dʏ�n�wu���ջ򺾵���%ؿva��6p��6\91K؀|�(A�G���^�萕�0�_���n�Gļ������O�J8��]ڎ*�Ĵ���m�y0��]@,db��ŪA�f��?�N�t�|���憈��LQj���gt�8 ^)�Q��4I����h\Ř�z����֔0n$��]FW����G����j���ln�Ƒ��ռVD�ĥSo��t�O��N���SB�c�{gL�5��Q�<\\��OBge);�B~��r�1��g��.��C9����ntx(�b[/���Z�]���R���]���m:N�TY�'��=e��FԾ��UK_��>S�Hy������pj��������V+Z �+Q��j❈6�&��v�t�v1��'a9�F"Z/�QG�L�������,(��%,.|��n�gT���;`��z²#j3u՘_bz~�^i)���n����aL��?�&�R�
X���t�.lg|f3 �y!�3Nz�����^��XJ�v��+���TC�k����3�(�B�}:�?�Ȯ׮�/�D.R���U<�Q���m�^ÏrF���͍�>Ʌ�ZK��qA�*����m�>�݊/���`���Z������0��r4z#����y�DˀS�V+$g&~>'����YHB�e��[��I��B!Ia04?+�oj�ׄ���8rK���qb3��hLV�{	Q)��p)��@%�BOt>t@i�&��1�,ݔ�z� '(���ˉ� 伺f�U*�ǩ�XD�^��6�_��x��5~w�Fu�,��D��	q�,�$�1�c�!C�RV�0��dR$8�{��$R��o��y�Q��;-�����x�*��+���υ�m��`D^�%˕�`��:�a����hh-!m��_��������J%W (�a-�N+M�uF�e�DkC���U���j[ԝL�<�cGR�����F����?�FHA�W��� ���Iz:�	��� ��`Ƅ�Ԗ˂W��{��|���[(=�VL��������gB�!Js�`-�l�wKݖ��R���{Ęz4�"�Ɉk,]��k���1�ݱ�Av� ��|���s'�%�`�F���O��G�����e^�Y^&�*G���`Q���إ�b�DH2�����q�0�c��8���HT4$_D�Ɂ���{/���el ���臤P� ��iPġJ��VQ�~��o�~9Nɵ_G��h�t�o�qi_ҍsۦl����5ʪ>��:�n)�}e����K�� *3^{���Ç\��k
���秴��wT���Д2IG��<4����Q���3�� �����	��)K ��WfIy?~d4�+�&��yn�-��{���&�S}bsk�GEו
a&a�.':��ĐWP��M�Yt7;m�EA�F��P���,�t[-��ĵb��oH�z�#!nw������'���Q��{e�|�Z���_�X��i���Y�z��Q4�C���9c*v��Yp��Q�����������8�=99d*�NX)�Z��F�4�S;X���}��a8|�l �14~���3N*J=�tF�WlX�����'[/.��>��lMЎg�����]��FCF~`Ѓ�E|��@|����D��&��yG�a#b߄�ށ`N?V�k����9�	T���k'���0�ܶ�Y�	V����'6o��?��@;3;~7�V���%c���$v�w��9T!P���;v���0 �[�B��J�&����%�3�:*���{�A}�Rr(g�K7J�ѮG1ϊ|���'\*��z��e٦�^q��X��7U���dh��*ɝ�ۼ����KX��`�