XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��cV�"�x����!-0�(/����O�v����DJ0�H��p�A�`jW��f֐�zU�_��#���\AV�v���z������������ҋ��
��+v��d]�4��^>��@��gVdu�
�&}�:`:r�����F��B$Q!��bٝl!����̥��!;K����St�� /�o�EI�:r�����c{�	�g+�a~	 á!p�(T�QQ:�.8 {�#��*���j�i� .��/�U؝�gp�!os'�A`�q86a�?��.��(��2��[��2� �]����������\�̣�H	\k{݂����1���!8D�d��Z��:#X��S������p�.u@�ٳ����H6�Ǣ�s��/瀩�a�S�O�0�s/9v#h9L��z�r�.�%��8 o�ЌD,/I��"��A��e�R��������
X�1W�ކ�S��>�)����`}��Z��W��@e��3#����9g����V�R�z���ӎ��!m�)�sڑ�	��#�}Q���_�����~kҔh7a2��n`c�=ʠ��!X����$?n#�n�>�v��k?�2��������w��ʁ�����H<=4���(�Z�z�ʷ@V���F5�lEb�օ$���=��ﭟӹ �^4eQ״@�L�5=���1�7t����ltI2�:�k��yb��n	m�A�Bn����<ٶq�q����{�`SMH�V�W9�7��j7���e�:&+�	��i��Z��XlxVHYEB    23aa     6e0QM���0"������T��{���=��D�ͻ�������'�Yz����F`V�HÐ�s$�����p^����u�8f �'Οu�x�(χ*b�*}\�X���ԊY�"����d�Cz��y7;lE���j�b&X��4��	�?��?����h]�_��F	)�F>u��/�jm�5�uKm��q���-Z�<ɁnxM�=/���3SH�l����`��ZKF1}�û& ��O���cWɺ.�~�x����w:�)2�t�F��P�ۥ#Q�[��C���.�n�o�_�u����:�@T:s�@Ct ��dq����DN��K��Z�n�/岕��݀�+%.�
�7�߲Mmp��p�$����Dw��!@<��0n�I�e�/��w$�`�6&��*�*j�aZݵ���Y�f8�\�8beA����(RFZN<.n~In�L���A�ݡ��,ͬE�����wa���ƶ R��h�R��<�7��g����;CW�Bb�j����2<�����J.����C�P"��"W}��vdt�GJ�K2�9K��$i���,�79�P��r��/<ޘ�:;��t|�nUIY9�'�_v�POI�����*�n���^��qknW�.k30,Cԏ��!�!�BxG&�7�P0s�H�4Ξ�;�D�c�D���֡/���=p� �{gV��$��a!'�SQ��H#�x���ڳh��r�2`f��?��F[(!k8?3���gu��o��M]��W�U`H����?�#� �@)T�m!���ڇ��1�xP+�jƋ��L��ߏ|[�:ȹe�Afa%�D�l٬P?��j�{�ל�sb띐ʾQ�ɾS��y����3aN5Q#�}�ꠧG2�1ݭ�Ia�+��:���:�;���nkzH���&|��>0U��K��6i�rp��SF��de�a0��V� 7"��:�ϱ3��w�N�jAXA�,�� �*)Y�@Q�?s�#�O*$�e�̂����ˋ���c�5�"�;d@�b�%X�����?��D���>m-;�>�����!��V^�n���7����3��䬠pgy��U����<�eU��-�кx�28+�1��Gf;?Y D�ӹ�ɹ,,�zor@. ��!ř�c��A_�U/�@�j�M��GjɆ�ǵ�<�ҫV�����2�_O����S�������*v��B&�j��}ӟ�� F�\���k�	m�.��᫺����H�z�]�bO�10�Û��sL��C��:�l��䋒V�C(��2�%��uK����==kh2GH�Qg'�������գDk���ښ�K��E�H͘�٦�p'�
\�Y`�9�'>���6�Q�w�mk�$��D��6����
�b�g�D��xC�${�x���a��qgZ����'��+��;�ex�Y`��c���.ع��H�c]b��&� |�!Yꄁ�A�š��(������C[�{����E#�p'8���k��آGz����O$���H%}L�?��5%7�U:�ݣ�ϞzL�ypֲ���>�O�~b���t?����)��뺁'��ƞ�!���
Ξ�����o�2,��I����ln�����Er�R��J�E�U�����L!����bilK� E��`����N��7>��?�~2֕���ǰFS�֘wF��y?i����7�-���e�b^Hr����
w��o�>A��sRr��x,�=�%KN���