XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���� 1)Z���vgHT��� �]9�!:��x{�X�	X'�xl%�����0�����9(��l���1�~��v�q�^ff���)��E"?�[a<���;���?8����cV��L�%�Z%���[:�2
:c;�9����z���<a�0�<��kY�zS�;���"�W�������5�*tPd0�����;�,�MsE �������Ƚ�}%�<o�l+"]�ψgM�<��ˣ"8�p��.�β�K9�c��H�*%���Dc�5׍k?�(h�� ����wژ���h�7��gQ���'� Τ:��,���iO9ݮ�7H�z��$M�"�-W�C.�nmk%�?|F)����31`��c$a5cZI}i���F�GZV�p��8������i�+N��3�p'73��5�Yre�Su|���=��oz#����>v1�䄛��"CϪȡW*kwPH-M=�� ���@.yս����H��&�j�[�%XB'��&آ	�m���h;�lU١�4,eO�:��"U��a�H�i�^���wy�$uH�C����=�����ȃ�[\��_�WG3��4��f#��4u�?����_�w�P�.'�J-�$>}�.�0Nȼ"����jBP�*>����L;v�j�(�����_?�A���Ԋ���}Э+J�_J�;��6����ܞ�!B2}g1W2X�'���ʌ�19��g��U�ò�:Pa�
򮰚�������S�	)V�n�����ƣ2�XlxVHYEB    7759    17904~Au*��N!��BB��	�����"��I%,����XްƬ��Vh;)o`K34\�h�(�EK�%JL;�ס��(R�r-GC��}?gt�3�*� ]�v�ӱ
#E��*��j�$�x�]$]��5��v��ܰY������6�a���YE !����3p�\��Ɍp�l��A��ӫ\��竄	��0������ie.pDT�_9����fq�x�$N��&9�MtCI��(^@��|�����t�t�*S��k�]��n�}-"YZDGP3Ǝh����͒�R`�9�}2�����Q�g�x}<!>��Sxhnpr��b��3V��|uck�Zp�e�P牼��.S�O�2���G�B��r�zs%���e�6>��J���Ւ�7	m�aI�6�;8"q��OA%X����y)`��mk���2�§	v��P~���i?��80"ҒO'��.�w�ar������p
�e���<~IMV�4JZ��V��uDf�9����io��$������M��(�_l�+�H�x�ƣazJ7�ɣ"�b���CP;O��<ҪK�"�oӻ��t�X,No����N�:�F&����L��[p�㖂f�w���->FظM����4�eª�d���2d �
UK����&�n��E
Ͻ���%�B���E"��w���H-(�ӌ���}�S�x����L���w��"���X�wY��ˈƝ*ug���l �|!��!�	��qם)䍭�S��__Ȣc���#-o%�����k��⌲?Β�;e�H�֗`J9�
~(9lRTݹ8�7�b�?�8E$t���=G���w�`�h#�.�l�.-�l�2��d�W����)/A���	�\�� ���k�r�"��:��F(sk�㷟�P\m���r]m��Hbx��˷q�EG�<qqRuh���=��6�g�'�pdWM��5�MH�2��e�t��y�ኃ�e��u:�~�0?�'�?�7g|Rsu<����:j�W/��(��s��sNg7���,���h#?q
֮��=�%�'A���r(>Rb�h��suS$(�<{_��Ne��>�{��u嫰�]�Ҙ9�EQ�/�D.6�x��5���Ւ8G���G�=D�J��������Z϶NV������������2�y�\/����()�/����K��|��=��^BۏWG�Ȑӡ�t���R3i�Bj���NtGu�o��M�RGy���G{1_[��W+-�r	�f ��w2���E�a,4Be��=��79�ī��v��+\ˠ�P�/|���ЊµJ�%�"�B�V�H�̜Ծ]�(����p��k��^-А��4�nA�>��%~��mj(`
�Ȣ�t�ѝ=���C�\}�%��J)'
���G��ٖ{[����>_��7�e@j�]��})���=yo��6%!����N��w�8&��������)�X��d�3j�n�+���ި�!NI��>�ދ�5L��(5��iI��c]�WJ0��D��e���Z��X'8�_ߒ$�
��=�{��U�Mhi�u�]TW�g������@���#����&������ު�WF$g���4"��T��`��+ 焰?��n�����p�&�J��E�=�u� �=v.>h��H-����+�I��K �:m�喩��M��@j�ȣ�L���@��H!�n&�.Ω��'n���|�J��ٜ����RJ��#��Eت|�P��4��] �sO4�P�;��wk�W�"oG%9���Մ����8��OƾӏL�Л�t&��cXP=���Z�k���L����#�/ruc�nGB����v�3a3�^��J�p�8��~�"��{�Ka&�j�"tܶ_t�%`�9[��&D&4yd����� V��C�j�3X����uz�H� 	�E4 %݇|[���Z4����2�	�0��
~C�	5�SW��swt.�<��L5�7-�|B����]l��d���X� r��K��֓�{�T9�Y�f���(�C���x�!�����+�pF揬7�� ��V����3n�I��=E��7�"��50��qa�U�S2U���Tw�-X���={�q���$2;��]I��%2�����læP�7���N�g�&*���G��D�{q�g�Z-�Ѩɿ��$*(�����6��sD�[0�U<��~e��1X�c�ܐ���w��N� ��a�`잕��:��Y��.����!�%��)Ȟw������0�,��˱	���Ȩz���p<��g,�<�\m5�*�/uIuO5�� 8ɉԡ�,�G�88��,\����c�G��$$��6d�=]��`fW:��_.#�+�t�u�s� �p���U��3��a�^d���q�8V�~�F˹�{��� �Z�9ԭ�Do��9�E�Z��k�>S��*�'���Z��{W�g ��9^U!-^ �z1�J�7�k��f �id��ԧj�%N�Z�Ѓ��D��|~A]nw�[y�g�ɔ�*>`@l���Dx�vj=��q	Q[{�pW��v3��mέro���'S'�W�+D�$�k��ȸR���+e�D�4��z�R��^�\���Y"���i��;�!*I͐���H�}Т�hz�	�;��rk�"�����)�k�3�I����t#�'=��A�'?�(m��4�m.Y�JV�b.)� ��x�d����\9 :�cy��x+$���xHܿ�D��%	\�hI�ç�=U]ҟ~~�<B�E�v�b�2&�̞9�:0M놭��@�ש�"�!�d\}a�j�cT�+9bG	�m#�5%>)��}���mŔ^�P�|��=��1觃�]G�h�0Di�3����Ж����/f�(~Y9�F����OA\c�Q�[��f�E�
���G�����F`d�r�j��������d� ��ڂu�?3q��|�]����J�����ޣ�D`%���sϹ����'+`���Bb�f��3w����	=������,xx��zkL���M�kf����_ 9d�a�{Q�l�V�Y���V&[�M1�W�j��� *%zG�yN�q��v�=P�݇ڸb���\����*���"��i7ug=ɵR���H���16�Z� ��/��A,ށq�+�TK�P6�z]8�j��)�ۤ��nI"eB1�B�����C4z�O�g�]C����\o\u�w%?@�5��-���4�ݫ�a�u������촣�ǒ�댁�b���0��G)dH����t}��+�P�;i��и��b(��dt�ϑ��.j�$� ��C�A0eTx��n���FE�}k�;�qSҿ� ��tM���UJ(�4}ġ���fȊ��_��,�_�o���7�	��i���%�KC��(�ڋ9��.�'	$���h]-,���� �� �P3@~��Q�]8G�k/�"�D���h�������7�q\@�K:#��	��c�\�x�
�W����ilC���]����_���]�Wz�gs���F��L.B����<�=�1�A�V�$4���
�(��O:3�I�K�f5��o�#g�L6�\���3�f����RJ[�%�wH3T�0I�<�C3b���y~)}���,<��$;y��Du~�F8��G���͎CD��;�Wh�(D �0��4c�����2��9�b^]�Rם����[���3�p���mA���|oXA<�ٕ��$��qѦzA�~�=�k�`��rޥeި�����}��J�B3�\ٖ����� �t_��9�*#�5�k��J��^	8�_���Ԫn�Ky��؀oGg�b�Oj<iM]��a�ǩ�`��:��U�Rxz<��pS����&��u{@�Z�BCi����#�����6JɪY�i����zq�c{p2���*cK�����(�1�,\��o<xe�ۃ�]����E��84V�{��I�wN��]�4�$'�E*���s�1��^�z������@����3(���D������p���j�[�Y|�;���!�|���Ak��rC'=>��Yo���]��=�)���e�:@E�h�;D�R�rq���t*�z�N�.�����ޭӳ�7P��6a�B毟-���?�A��UܕKV�8���<eK�F6<a=i����70m�oO�czy��,!KzQ��1`٦W�e��lil@mz���I��" ���IOi(�@P�SB��s͍�R_t�5>Oa#).n�YS���sS��ѣ��Lzٷ�6��R<ĭroH�!�b�҆�+>*�bј�,���Q�vʃ���䬧TbmI>Bs��L�f�LKJ�~�D�zҿ^0��$�v�����&sXu|~V_1����<T�u�N�qR�l�)O%��b/d ���l�)N��t���w�AAjW��Ԡ�6j�Fs*~?,�=pzDK7�@v3�E�YgE�^yWYS�1`f6%���mZ>�b-�64�C˄������H���<{4�H'���ץ�mW�+��d'gu��PVN��%#�v��a�,�/	�]2�'�>����Et4���w��d��(P���*-eE�?iA"��nK��$��+������4�Ю؜��js^H��y�6ve�_?�����蔉�L���t���g����TwL�*s���f�:���#r��Pe���>(��:$Q4������x9
����u���=9�n˖g8���aC���$��.�!k)�L��
g�c�Be���0��m�+J�jKnU�l���@l$3�ɜ�:��K�����s��$	�ڦ�/����{q�`�ۚ�K��5��L�ž�Z���"�a�f������8J`Q�ـ�L�g���{A���Hi;�BihMk�xb?�N[�����^�F���h�#G���Ep�ņ�O�x�Oj�Ϥ��?�6ꤪHcʈN AyS)����X/��R@���o�fֺb"�ֶ���霏�ǭ�CŻ����y��PoG���xy�-��Q��,'J�#��Nx�bԴ$,�G7.WW��a!��+�"Ү������kO��7A���c{^����Z��%�X�v�7�6�l���O*I�u;�j�1^Gk}�~��'���"����V���F=xb�Y(w�r�fm���y��E�����\� 	?woT}׿��	��/ɏ<ym��DO�$+�Ѿm)I�ܧl�I+�,'���>�y�ہ`Q�������ϝ��s?m��m�ii	��&��-��A?��R�b��O?ɨ��KoEV!I=�u�Z>4f�3���K�+�ZRu��9��<��1�SƼ��4���(�V7��Pm��!&Ib��v)�E+H5�:�^Q9;��_�Y�Q�S,�@��eɉ'iuZ�"�����.w2�9-���	 �j0��y���s���	�wzTkZ���V�Ul�_o^'S��7�KzHr�鈟��H]��Fb6�G����6����
��9�����а��Ӕ��|�%�{׌��y�+�u������z�t���	a.��ɳ����sG\R�_�-s+�w'�&_�Lx��I;�+�vTZV�^�$I�*�^x�/�T��7���X4�h�������T7Z��׿����9���;��L�QY�so<�@B��qي6�`5���2�-:���bx`f��>T2Pey���_P�6�k��,�����Uf�{ձ�B�M?s3�U�Z>W o�J޲We[�$E�>�%3\a�bP�����ݙ���O�2E���{c��{g��^ވ�.?=Z�����Q6��
^��l�^�Š���:��1�qv�{n�ޚ���mŊ��:��ӈ�� @���{����J��[jW��\{�b�W	Xh	�����Ok/���h�]���k��W(B[���� ������\�����2�C��K��^�g&x�0��������{*������yv�l���H���)8�i;�h�~��*���2V�N�G���u;���<2�����M|�����J��e7{����