XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*ڼ��ZmKmY��([�򷲩�ѿ03��]�!�x�o�G�.c�����5����Ա�(������+X�fh�8{T�����X[u:Yh���y�Y���9n���i��h%x8����ĵ�Mr}:1����̍h~*�-9����n��%��e�ގ֨dq�n�ė�\I��Bg�WfOW��њ��(�ˢ�~��q���GK��L Ņc9WͶ�v�w�#��,x��.�胻�_�8�����6��S�#Cw5�0ck�=�6�����v͟k)e+��[WW��]ݪ�A�Y�"Z�Å�}�=I��c �!�$Z���1����l�z �6�=���!�_�zZغբ��4�,���>^!���=V���F��P��n�SQ�ͱ�{$�ә��mM���������6s�Y�oP�]�v��.�SV��:�P-3sN=�^��w*�ځ2@��-�g5�F L�<F0���=�YrTs��'��]���tr��!M�Q�)f2�uJl�ܽo~ˆ~�t0:���oM���6�A}p�pʷ��'C0W?�ɰ��BP ojW,`y��L�|kl��`�\�����beLu�Z`;�}%m�mC���;�%
�w��A$*�Gw �4@�x��{1n`�Lu�v�\����*�w�P�t"�F����-�����O������� WXO3�5� �#+�_~Ku��+�ɤz֌��gX�jP�']��j�e�g��Z925��H���j�u��6�2ޚ��9C$���2XlxVHYEB    409e     e50�3P��)��hhP���0��Oc%�h
���q��}_�"�S?؊
����v�7x��Aj�������I�����T��}���_���8ˇA��jwG����D*���=�!�Ȍ(3�;��>��ئ�jg)�D���Q�X�t����r�.�Ju̡��ى�
��&�C���*T����;��
z��fx�/~�N`4�!�[+��|��>��+�cD���y�[/�+���N>g����(tcN�S�U��u��,I2�BX�&�}h���mX��KB�fh�  =ITꄐ�[:�l�z
����"��[瘨h`��_6\�$!w�r�w�D�p#��%�i=��^���7
�߾�.�u�H�Q(�A��2���� ���7kO�0�j�b����mʸN��?��or��nQ����i�7_3u��ל�W��XrWi��+��/=��w�^7yBdt[X�+"��~�O�s�O��l.�9����OoMt���ʶq:�"{vYW����?�<qG(����=�����;�'T� 	w9iL³I��K��%L��"+�S~x��9'���nqz�~�!��i�T��`cb���sޞ(���s��s�6�j�4
Z�nw��� ���XZ�Nki�6�ӿY;Y��P��9�99���%���47�n
9��~���D��ܒz�vF�$hb�����L��\�3FWd�EyDk�}w��4s�st-hn�' ݺ�*��\�m�q�̒�g�+�U�0G�#�1��6�A�BZ	ؙ�x����*��S
�{&e��1at�&w2 t=��\�\���a���e�w�0�ע�����F7�±�n�Qdk�m�h2�D��^��x�y�`�����4��y�YU��`Y@�G� =`�	g�I��J�3���Vi��Kqw��a\��GJΟ+��C��c-H�^�*�}Jr�+�غ��j}~������ڳ�Y��3���$�>*�u�	{h@F���@<�Ma�H��P�+�Y�����'*D�^��Z�F�<�Coc�Ǘu A3������#�5�nqx�K0F�$;{���^�T��5�i��R��x��,�/���R��ٚUguVGLpp����G��Oefq���j��4�4�EKd�fm���YCq�u�]��p��@]����H�+�p�X�Xq���'e�`��;Y��n8�S��B˚��:�u?��.��RƘ39�E!`����ݓ�tb��%4���K1�4�)[]��u�P�*N:N��B<�0���u��=���dҟ��0�o`���J�R �[`�nB��q�
�������5*�!����O�:�bX�~u>�������dSS
12.U{|�d�h�b7cC%�.ITC:0�#� L���\���hI�{��D���KU�vz
��|@��
�T�$F�6��#��un�)� 2N� F�,b,��)&��n�Ft���2��_���IR}��j�	l%�E2,�i$1)��Qg �~Y��VRe����=�����;�R�{��؃z�I}��-w�z�9s_�W���HViD* �UnVPt�-��9lB�
�.��\��/� ;��cq+���*���Ec��E�x�`���0���9�
���p���<+�|3gJ+%i�����@n`4��O���px�?@앧Oq�T!��2+jA���e'У���ABf׋m�4"���H�o�8�s��f����݈����*��8)�#z��w�^����+ů25qP������RV�%A|���9��O��=Ù���<0�=�W��n��ok7��?�`���N��(�_����!��{��7�g��'�Xl��=foB��TB�K�X�^l�$���D��΄��N�?��6,���
]6�CD Ѩ��$=D��SYE*i�����aS�vX0!�V956qX��F�7���:�<gw��Bd�<�`4�[̀���h��2>��|��`�x�@��A�Q/�>lx�?��-� ���g�R�GUa�<���N��x~˝Fð�]De��b�������IK�P?n��Av��VP���Nk`�Gz��C����1�]t�~��#���P�a��:�ߠq>R�����o�s���دB�+4�!�"�XD����Ę�Fdb#9_w�G���I-%�޽�7X�~o9$��J��X�G��֢j� a�I��E��IC�5u�i�kɳL���bĤl�7_���,;е��Uܨ,m����,ԗ��#�f���[ J^�laK��"1��G�6b��9��T�1��p���f-e���N�-A~�A�ʡM��Dk�}����"w��b	�#K�g��y؝ɱ�4�A�?�㖖-.�
6ɉa�f�o�{�e�Wq2��W�]i�$"gН3�5�a3MU\�iO�>��O����_�� �� �<��c�gao�%�q��-���4�E���x!�N�8�r�a3�fN�B�)��=�T6�<��%�w��oIbz��~�w
� �ܐz��&-km���B�U,�Ⱥ���܁'�s{&�-�w=�tRfD���q������?Q��S:��,���*��[Ԧ}g���������5+�؅�-�*�SBBpN��a�S���H�,��3��%���I[�?��������V��� m@.�U���߿7������`R ��w�P;\鮒 �,����6.^O�/-~w�Ԧ!����ƴ
���:�\���RJ)h^;�{������k�"\�)�'�-.S����.��]<b*�4K��Ȝ��Jg��wՌ�@o\�X��5�O?1���;`�^�sE#d�H�+�q<e��/t�"]]p����g��������KU�6Wi��q9��S�+}�`?f͝}i;z)�@�<��2� �;��&�.x|�m�&;AP���X�9��2��P� N�ܮ��L��,����pnՊAa��J�-Ľ��?G�j(|�J�����Ǭ���cs�@5�I�r�.����N���ӳ�oUڴ.YTz=�a�uD�ŸF� WX�q}d>R�iI������Kْ��W�&\X�Z�v�+��V:���޲��U��Z��� ��k�j=�-�,o�$4��^^��n�ºǠ� �`���ઃ�4�4���-Fb�YJ	x4���Z��B��9��������0LU�΅�?+6����[˙������g*��<ssD�(6rZQU�d��w����_z��]	x�LK��y��-r&)�''�*��R�/�r�m`��Q�V�C�6{�0�Jk"ў֎,�7rG+pr,�p���]���i㗎�cxX�x)�h��A9�Ȳ0��"�5�\-���w>vv��BfKm���{<�#<{��2�^���99�T+�牰����^��1]q��'2����>����0�.Jɷ;P,f�ڍ<0{c��R��
;fP���z��{�e�J\v���j�{xD��f�S�:躟%�(�pU�ǥ�\<얄o��FTZ��m~4|r�2��	�D����Q�����E��]�B=Qu�>L�A@Ma�3��v��E����9�K����B��ɸ�_+E�����y�'��y��rM�%1��K��0`!O�xo,˪��aQc��4��-�BE��NJ��;3V������5 p�үF����t��