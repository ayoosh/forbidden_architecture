XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Q�R��Z��m�e{�:�p0PM�����ƫVynx� ���˥�܌�s�������PXw�`��
ṯ9������GB��*pB�f��k�/�7zG� �'~�j�{� ���6<_������쏊�V������)�\���xz�4���xS��7*��v<�ʪaк?���->^���~�]��F��c���z���I<��Xǥ6 ��!�-0k�H�mj�(քL|��A�<k��gȪ��#�+Z�\���bsA٧2��Z�0������y��bpU������Zl�DE=Ҡ��]�Z�!�l�<s�N�;�)�����*��&�|C+O>Y%�6*���&��
X%�)e��ay�LU-��k����&:4�Y<���B�7X�\ǱLl+�`EɒE�*er�HrD�p�!��K�ׅ9�{}b$p���{4a^A�?�V�)9�AyEڶN�]c ���y���o�"+nuw��<;6[_zcO�m.�T[K!D�'�$@`԰:M�2P����0r�恪���Qv�r)zUR�4`�!*����w�B��a�yQ���uJ��R�q	�@\=Rd��f���X�v�n���yb�oM;JR�'L)���1.��>�Op�iJ�C(���ݍ�k��f��r�<�H��49���C�9�os�!,
%,%t�y���͹��y1���K�:�е$�5mh t�7K��-ǭ�_��8״	�.zS�@���nw)��s:nD���j0�.��gXlxVHYEB    aa46    1e50��Y�� q�	�˪DC�!տƣ`��6W��v��J@�Z5K�'d�
=���ܪZ��x^}x���m�8�%�e �\���1jtwh�!R0'Ǎ�eKc��W����Ө�*��(����ܗ�hI�g+��QFiE���t�n�,`a�z9H]ܛ��w ��ݯ��S,���sD��`�a�y$�?���8�1���8gP��ҙ��x6J�	�|���(S�&\��~��AA	R��xJ�W/֏�[A+�[=��۱<�}�wק��VV�@ls��N�l�sl�M�2��/�~�'+eH���h�w(K|�qB� �f*5(p-�ϼ�f���.`�h�>�t��#�����.G;h�0���>�LA_�|�@��L����V2�<�,Û�4Ꮂ����b����G��bu�A/��C�5ɑn^�������믾�@c57����8N�1*��o��~De6/h�e$B;ʲ��\Æ�x�]���!��F�3r�lZ�{ؿw�`LZ��_׫��r	,E#{6���"B|��f�@Җ�PP (v�@�Gb"1C'�8YtC!���i鮠D]�'J��O>�{�
h��W7��Aw�w��f�e�=4~a�;'J+�8����M�Q���z:�˗�4����W��Nk�t�����,�D�}@�t(6��S�������$��mn6U8>稌��T
�6�3^�`e�1�r��=��͉��&���zY�@"��ݸ���f��qs�\?�M-(XiM���,��m�q��U>i޽oȂ�/ɸ��V%���b����J�5�����&H}�+�=+����<��
G��U����i5B�vzT���L8]~o�Y��$Kð淠�k�t&�y��`7���-f&u�lA(�EŁ�[���t_K<�Ey"h�-?}{�h�P��C� ��Ǵ�hG�T2�d�ʯU�2���Vb��y@��j�5^�Y
�����= ��h�>���(V�Y���$��^�̎���f f23[35��{8'�3��x|W�&(�Y��07��1�@ƿ궵h��8���Zr���?��'O�tɤCw��=K,)�"�gۚ��I�pI�vݨs����I���|�ǜO��X�4[��,�O�;����81�1�$��K��M���V�&y��1P�}��F��T`��}��}% ��u��^H���RA���/�J:gn�l��8;���+�M�E�j�$�Ņ�t#�ؿ-2�L
���dV�J�\��c��3R�f�z|d#	����7B��P.a[D��h��`��C��v�EB��Y��F^+�P7�	T�p��Q��EN�X�X�7��찬�h�rK��ffѾ�7͈�o���U�C8���;4�-7�-�)ܔ�zb�uA����e�Qb���L�%�U�mV�Kֹ㬮k_�}K�?�M3I�Ǜf�;F�ટ��%R��S�)l�q��$p���>������ur�e���b�o��R�CS�-m��`�8��d?���P-��9�E�E2�Æ_(�E(��'�v(�,ޜ�$�|A��0�HO1h���Y����3z~�X�0�A����Ɖ�;��!P%k�^����S�g�F}���
�\D~,����2��{F�:s315��ҫ��e0�ul7�5LtpB�b��dQ�W��r�� ��v�zIN?4��Z�{_A��\0��
������X8x~X6	��p��k�����k��#"�E�߆{�����H���yg�x8f�A��0(:�J�\�C(���P�H�*��2��`��F�isjE@M���=;ad3��H3�OդM._�a����P�nBPӈ$�<��7 YD2٢H�j(���Q>�����$�$��S�3n�a�m�r,a��`0N��^��y����S����%�f�<��wv���oDk�nJj�7Zi�`�+�y� �����"C�-��&��ޤ�\���4)�5'�������@xo
�gUM�{M�T��fs��N��QrDC�S�_"�|��҈��>�(��z�GM�H�H��J�J�
�s�G�[�r�}�3|�!j탉��<'�~p��E��Gb�V�{Y�Ж\���g�yB@�g��v.s�ǎcD�4bKZˢ�O��`��4�p����6��5V�~�?u��������讦n���PV�h����KC�߁�%	��\9!]��	�@R����۷��H�ޓ� Oz�z_�} ���1��2�c��~/ο�Vvl��ǎH'a7^_�J}�+�y���$��uA#Yqڛ���p>X m8�]�7!��4u�ĸh�����7�5�.��焋b�[4c?�x��1E�"A6H���aPL�-��A�g�{IT���;��I����fO�R���9gFXF}�f��)$~��w O�v�K�� �b�
�� (+�gT����6����$���.�u�^Qg��.��tU͈ ���d���w�Js]1��y�$���hoӑ#]l�7w�vG*މ�O�4��I3�z�;^���`�F�.�Wu��� ������=�������ȣ\L��yi�P�dߏg��^x��+�RyR_��kτZ1��aa�5�Eu(F�pz��2�:_�7���H�47��wK�Xq�_b����A�@�����|q������_��c�̤&����X+�eg^�x�^�2�
��*�f�@Z��s�EA-mv�}��P�T�9Kn�h�¹��t�<�8�����F�wL���Z$� P�?�1����?���γ�G�_>/���b��0����r�;�����9�g5ɂ�:���s�M��Yu9U�qC:>J�[!�h2�Zk�A�.d3��7���|`�w�����N�%J=ʈ�W/�p��2��:^�i���MS~�.k�YqX��l��Dѝ�3���Ӟ�|������v�Jsl7�2%��$R3wlح�/���w��OM�.<d4�V�����6D�}���Ԩ�y�/ߴ0[��^��Z�]&���񤄕T��A�2��9Gd���S�+/�-�F0����M��X�$��W�9�N����V������Ʈ@`XgA�*o~�Z��u+�=A�Y�����UT��c�!`8�>�JB�W�l@Vה�c���N����"���Sz	�&9ZF�4+�3 ���5ي�Q5%�M�Xs�#���EvL���-����X�5v"(/G-��uړR�`�^I<�q�9ٌo:/�Tw{!�4�9?�:Zs�DL�G5���P<n����M�/�60��u"+݅�NM�H�k����|�����,忆�u�R�8���`sń:�>i���0����3�nD���r��7�_�H���K��.��^A|���ױC�&�¡,�c�PS�dҘ	�C����j?1C��L�Wb�Ͷ
�Y��Q/I����S!ȑ�x�wi��'��O�6y�!�k��8��n���|lO:�_��|E\F�lM�J����.�\���.9�B���D����s�|����_��D��%l)��R����0'�?!�=+si�T�l�wv�$q�����|׼���J�T.R��"Mai&�j�Q�Ԩ��{`*�ߜ��)�59v��¹���N�&��1B�۱!��M�,E-\:������8}��s�i�A{Ƌɒ����tA����Z�\�v(bWt-��8(��9�q�mP�`������/�Q���)�B�2��w=| �aAƣ�U}�-ᜌ��@9ˍt��O-�&����hh�U�逥�o;[ۮ#}D;�`�4.6
h��C���dq2�<Y����Z��˔и�:��[D�-71'ΪJ]0�͎�����m�V9�`��즫��M#�!�ҡ!�{����%��������8{���x���5���o>���@?|_t�r#|�ѭ�~�3�Pqʭ��KP��4Io&\�RE��"/�ߦ��@$C�j1)����Y[�Qnْ _��o�6�-*35��fyoirE�uv�A�5��_`R?<;KC�B>��ׄ�k����x5��f��� ��c��M�1Z/ ��,y��(5�[t��qu���XO��]��\~�F�_ф���kk@&�adF��(�B��EI��.��J�����à�b��
.������S�0cb�h]�������'G����q������m�%��-ʱ�B�$���=�)�晍���1)�k�:D6br��Yl;p���w rUv�BS߰l���Em�`ܧ�4�u�����M�I��m�7�l�zQj� 0h|�E5��+���=�M?�X�i�2�V�Ye#��X�LB����Q����A��ˡ3�4tn�=���vZ��:�2A�.��Vp,�RE:@��?`R6��<MyK��0����${��ϛ�ܥB�2~���Y�P:6�@[�/!������`�����S����5�q�<͸�J�.����ד�����"��(a���' �Ԓ���Y*Q��Ꜿ%��b���cm��E��@��0/���-��������-
���l�*�4 ��ȑ�� �7/�A$��g���e!a�bn�S�C��_�/v���l�{�+rq���P�hS�O�Zw�d	�?ZQ��Ƙ�s{Io�s�=$�(�9p�H�ߞp��~6{�,��@�&؊��78��L��=�t�"��6t�{N����B����j���l������X(�_���XSBl{��d P��kK���_ѐ��/�]g;��)�>�bk[3o��[{:�x"�Nr��G�T�N�%�Bb;~�2�q\]��HiSsU�����Q��8���B��:
����G�c��@>�1s�e!��8��XUMҪ��Z����>W����,���.�I���T���������I7{!d�E|C����,��6H&��<��(Oٕ*�!jDHx��ɴ���V!��׭H��z���q/`�%��J�'4�0��}�6&���1]��� e���$��M�IN_�Ч����T	_.�XБ�������.�۟���`�[�!`��{߹�PP�����38]�Т��E��#�? XbX<��'�� ��>�SȨ@���o}��<�� �Yʒb�[)�o7W��~I��7���B��iԅYcA9���6���gZ�j���ۤzf\9)&��bq��d����i7AoExKj8V��A4�Ƣ^�f�WkaT�p�M�	���^�K�<��:�P�ƍ�'?S��1d�d�k,�OIX�!?�e�9EYI���B'�I�nR�&��?�*���z���q�=��& �v���]�~d�Ԙ\��w�Ȳm�c�^cX�9�Yg��^$��V��F��GU$R�.LOB3����B���n���o�X��D�v���J3�O�W;��9%��ۈ��D��Nk�፶1P������b$6d�3��;ǖE�]��ե�ꪟTl��΄���E�u���\�9�Njs�����ٌ�α����9���,�A6���H�G��c�mz�6I��dfОb*g�܌S����_�]�r�S�8P �l~^rC��^i��l�h���Y;r��`cB�ɑ	?XPR��,������c?��F����I�`ߪV4���8�bU��@ȫͨ	�+���]ũ�Ъ �r��VŇ�(��Zj�:W�ék*���ؒ�Т��bDH/�8ZY����	�:��i�w�Qn� ��>��e����b���]���������������@�
/��|�`�����s ���m�NQIÙ�w_��O��
�3c�E�7��عXQk�G$� Xq&�~��3|(��_台����U�*��,���U���I��C8��qT^6|R���:�^c�	x����Utә[tf�:3FKAe?g��DSC�\t~"_��@k�q���6��\O^y��P(����"��ݾ���70e����������s�։@<
"!��)��K��Yopzg��uW���f�}��$�P���=z7c5��yMŦ]�g|3�@ߓp�\Y^c�M������@�y�_��`����m��?6�1��P��;�㍳�ݤ���Ӆ;g7*�F��5�Cv��L�rK��ȓZ�;$<Q����]X#� �����jԧR�i�_)/��Aķ�V�Yd�[�ވ�ס�偑j�3J+�߆l�x�͆�t���k�B>o�����?�~z�-٩��K�آF5J��x{?���={%:�z+Ǝon����*���׵v��"r��v��;��P�\Y�Z���?�f;�������E������N�<�އߺ�k��̿�g[�W�w��w��:�bS7�j�����z�&�늧Y�i�v$5y����A���O�}}U���V%��w�����s4$��!�M�����kQ.e���>4�F �پK�iB�P�-n�`��g����A-'�͞_xn<{{un�8� ��LM���]>PG��ec�j�|��&�Vu?��e�{˜����)�g^�u4M`��U�k���wAs	l��5%e*����t'����)�ה��ɝ���a߹O��ɫ�H��� tK(_Ǩ��wi��b��n�67�0�'��Ϧ&ꅟN3�I�wQ��gX�[qK���:�ޝK8�!�l@�l8`���[	��u|���"E�gM~��,�D$���7Ͼ3���?�O3���o渀���L��r��#�9��OUvD��<j����Lڳ�a%c��������+z�a4������gA�>P�Bsb��D�-{^S�{Ɋ��3
��Q��6�����������W��&uO���t!�m;����������u�(��f?�E�弧�>V��'s%�x�5K㖾���)����WQu�e���L�*�Jm9���ӓ����� �5$WZ����j�P^�kܚC�3��ZQ��
	t��v�4�f�k�{P�� ��]^�w�fH|��ű@��I�n�T�Z��������88ঊ�=@�ĥI5K0=@Rt������ֹML�b!s%==O�W6�^�2������
5Ic�Jk�F�H��6�g���a+e��@z(ǳ5�2S�����j���6�4B��]w"u����o�����^	�FE�@�&�N�. R]������{����ǀ @��i?Xs|*�ר$osT��}���ne�x�'W�m��Qs�,,R��Ϧix�i��i�U��g����/�����*��)Qy�4%L��5����#���l���#��oJߙOy����{[m�8r���"j'"��˭.Z��T�-!�z�\�ͭ����S�xʭk�]��|ӆ����<m���u��E�����ȵg�U�Ӟt�:�l�'���%��F���Wa���ߧ�w��.rK�*�QD�����h�?�T�LZފ�'	[�y�\=D"Oz>�$��RX���[�qC�?�B& ��zTFO��ELDϰ7b(ng��kn����,|���t��4�S����D���O,���ޙ�.dD2�ݰg9���"�����C�T����B��H��u���{,��������%���B�m�~�S��>�*Iv:
E���n:
��)v��$	���&"��"��`�@�R2�&�{#Y�EKr�7k�i�=]lD�����ؐ(����s��qG���?����r��pj�