XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=f����|'��!h·;���IF��tS'B��l�^"a&���m9�'�+aPF:JG���ɟ��]��KlS����;�'p��B�@�q�7���x��<���r�Z�M�!��|m�ؔ.itE�s����h�lDo�̵Lu�W��T�q��S�e���m?���^I=�q��!;ʍ��+���!���=3���n��V��B�q�[c'��v}�W0��.>��J�����_"������
b�-rz�-�����z��n���:E�
`��h��Ba: JJ02)�h_&'�L��2ȫ�K�	%\�S=��M="��m�`������FE��	]�b�i	]K#�{E�i�+	׀gJ-$�=k��E��'l�ay�#N��}:�X�*'�d�IBD���Q�p�ž,~�Ŭ�&qE׉-��L�!bm�=�>$�:�'P1?��fQ4R�[�|�,F;l^}1&�Yq���,@2F�$u�����Ur�����"�<��:g+F���G��֐K;�N�Aϛ�<;����Y׹�v~�g�$��-���:�/��u��A�`~��{)F�m���<���!vj��,�pE���b1$���'l޵$�Μ�vww�E]Ŷb��o��W����^���f�'7�
�e�*���b��d?��Z��O8A4�r�4/�EԛR rX���������v/�A�fh�p��ȰE�9�n��Q�%�<� �fdh�w�	_�mpea��8[��}�GPD�
��+���Z�
�
ԛ�����I~�XlxVHYEB    7744    1780@8�E6bm�q��c�,���Խ��ZWy��H��7��)�\�ͽ��jB��{���7)��������@1O7�]FкE
������F�Y��zg�@Q��"P�W��,����﫶��v�.�����Z|�������.�&�2�� Mi��x�ir$�mzZ�T���Oj<��Ӵ;$[2��F8�ԣI=$^<��j5B#��JL�G~k,��.�Q��w��Է�An����Ǐo"�$�6��=��E�lҪ%t��̦�ZO(���_��_�F�1J���?��a���Ph�G��F����'�ѡ�3>�����I��C/�J�����Q���3J�̽�aH�?8��N5����qAӽ�v��g3Qz�u��K6��xo���:Wm�?��<�׼7��W�b���-�[G�;�.4秖�PFޝ��X <P2��\0Q�_�WGR�|+���n�������_�����IC?"�V�����'=��&�䵞�@>�òf���%�oq��P���n�O�:7��*�����3�+���ǭvڳb���V����ʷ�v�!#&�T-�щ�+��$�6����"�d�ag�3:�C����9�r$����>M�b���o��Y,�Ҟ�H$�*�U��'�Mw�U�BpU�A<&;���ƞ�NexmR���@0���%�����u��e��%��ݫF�un�HVB�HJ�؏
Z/R-j��-�=Gj+K&Mˍ�����,�uTFq7/�:�ӷ����t��4o�@�L���6����E�gx},�:���c�U���"� �5�lr���P�̈́���~�,������������!v�*!7(l��iȚZL=_K�5j�A�#6�w�}�6,G�����im���Ì�cB�࠹��}W�ɹ�7iR�,��#sZ�4ʊKv d�cC|/����ӄ���pO,`���Zǜf�E6�R���9ԥ!PYwz���aȚ��R���WҶ�	Bh:c�!�~U	�t��|)_�����#����ׯ��4�%��x��8��Ǒ�Ƕe��q���F�����L�<I��(״�gk���t%��� nz�>��]���,۳XzZ�d��ӔN���U��U���0%�3t��vr%�F�bE�J6֩��j�N3win���3�b�h��E}Ҁ��#s&�'��R*LiC�ɨ�ڧ��b����AqZ2
U������7V���$)�^��>��/q"!tW�n��pS�Q�L2�7ճ+����s/sx�bWǔ/���I,q�?�u�%����"�y����G��0�Zw�W����&b/<�����M��`�&/��{�:���@5j�k������}�s���4�}F�b��/�\��l��..r� �('������W�8')�r�g�
V�dG�_q��f�ן72D[i��a��
C�S���lgn�a�䞘i8���^���c�c׮�˓,�����ZҪ$:�f��?��_#1��BO%q�:\^���v����`�:O5����ٞ�٬��GϨ��@��h���7ˠ������.�����[�$�b�o�5�i�{�|�9������}��;�Y4��kE,� ����q�!��9y�X=J>F��[�$��~�B
<�����Kҧ1�Ǫc��`���	"=��'�Xz;q;;�����I-�!��;IF�v��|ˡy;_�����uy�zNO{��zT�i��|�	����r� .V薁w�S-�e�A��p�t�]Xq+��-����h8k��6�������t{}�-�T��ycq���ZjK�e2+��C5�f��:��kR<ez0�����5鹞&�<H��c^^�d�]d@U�#��-�t �ך3L��p��@Ȑ���8�h!l�UNކ�F�y��6N5������"��&��)ǎ}���9\s�zi�>Y���
���(?껡���@fc��A����'/ݓ�9ك�w$hn�9"f�E}�7P	��I��3��@\#��p������5tY[C}���4�tp����j�r'��Y�u>Z9�=�Z�3&�5P�z�����*�w��
]���(�u�
�ZT�N�]à*��L����u�C��AC��~Uٮ%�G�b��^⬾��V���=��w����b�������e�����EZ\�Vf�;�������.�i�2�WTn�cb'c�����\g-z/,�����/\Ǳ�+�S��'Pũ�Իˠ�nxX'ڙ3�gW�m x+e��l�ʴ>49��G���`U}��-��W.���lv��Lk>lX��۠d�*���×��Ym0ߖ���r�I�r�	�NBڬг�p���e��8��d�F�;ZuI[s��yW^鴄U��V;ׄ�R��i�V�
�N�u��t�O�vOS����4j8L�iC�������∮}��FC\h�U�e��M�?�<>�k'b���Al.\�F�(����"�e)��V.Q]s\+���'�ewv@������N��3�-]'�>d���W\���~<����XJ�p\��Ap���d�������~A��?����Ǐ=/ s{,�V���yH+i�-�o���e��Ǳ��|��,����ׯX�e��f�.H�.��z�Tzx 闪Z�P�-���:~nb;n�Pb��	���dX�J�H��ڭ��-�墨 C��[j7bfr�5�J�OI��ќO�
�!(�áH�q�&�cc��i����/�7�[\�q�-�f�x����jA��גS�C^�� '8�Z��h�Ac���`���O�\ w7\����'�;�l�d&1�-,��EM��!�	�Z=�w�b9��*47���XT$�+�����<Ht������U릺"�}b"��� M
����lG76N!�����^�9�I�ظ����%��2��,�ބ��wfWo�x�l����檷�٠�L��L�G9�J���Iߔ�0�<�˽��UFKc��e_oƯ�թ�|/(��v��7��x�/����|���A�"��ܶ_���R1�F[�����I�+u�����4�r�^��ڽ���ϻ��1���oĿ�2I\G��*���߀�CꙜ'(s8������*�i��F�2���&v��J.Vz Z���]T��v>�(�|;1� ��꾴�R��~���8s��epaqQ�/��)/T!
vd\�s��1� �/��p�vX�p#A-��&�aɡ1��vr����V�xu[�6�56��,;l1�U�E�2�m��h�իհ�W4#��4�a�b�c �A����^�`�>7�O�k������LN�݄&�d #�T�漌u�'n1PԄ���ѣ��e�?�-ݛ�Gz�C��������9�&���\sA��wȧP.�Lj�̴n�aƠ��M:�<�D�yX.w���h,5�x}��*�Y�������x�K6�h�$H�F���α��?��%�O�.#��ho�+p�
V���@���ȷ���H���>c2s=�n_K�ƨAД����r3}L@�vq��{��+^��1���hu��z̱\$���E-.�TO�CLp'�p�&.*S_��7�(6�^� ��"��sʧ|S�k�Dh�%'���H%}˥ n�T��+ݎ�?2�V�!��KcDjA�s�d�1��^Lw(�wC���*��Ox,%�/�7��1Ck�\|/IN	��j��/YI��������~�F�1�j���KP��6��"&a�r:ts�	�E+�З7��j�[�U���XP�HC�t��<uK�N����	9�MG �.��p=�s�G�#��hZ�J���>��uf���s��+�B��X7��_0:&��u"4�5���J��C4}�u/5��>`��t�����/��apPC�l���p���������3�l|6+!�r�������k�_�Fv��]�Λ��rMu{5 ��S�t1,q���z���r��:��m+�%hGIG��{L�𲵫2��Z_d����yX��i\�i�aR~`S����������&ܞ�A��>�<�Cl�an �}3i��>]�B�=�cwF��mv��/��n�)!b2	I~�:�� e�L���y#�ː/5Dx�T��(�j�v"-�) <��P���S���Z���[��"-���{n���#״F�L�E��O+�=$Ytd���P�Ht�=��EX����6ה�@���X�3���c>�o�E>�x��>��͡�A��V�yu}�ߘ�f�}�+K�X��}�z���� ]
�o�
B��?�����nAR���;F�R-y�.%D�,�����S�8��YFN���j��n�]9k@p�F�H(�Z!�=�f���>)�*�V4GV	�Nu;�\�*\{�@m<���ӕ��	*1�T^a=���m+4��҄�ƹz-�F�^ :Do���$<T>������K�ӎ>z����N�5e�`5b,?��a�2���]�}�{�C=�>M���y5ب����]t���F�B����A�؀�$�	�v'E�:ǿM����=d�pr�v����{r��J�����)^���f��"k����u��cEa�>�W^����S5�.8L�Z���?- <�,�u9M(^�؊�tJ��N>ÒeI�x��,��		M剕XN��!�T�2�/�~��]M� s%��Cc��h�"�v����j�JK���m�|h�@�<KUE�P����z�e��K��".FA�?���m��.݄��JS�r2��\胶���X��-M�f��M>����ϋ��S��R�R��4NJL��3�
p���!�����̊�I��� y*������{3��Œ��
�C��Mh�]�N��2���X� ��;g|��4�ŎN ����]j*�`�A2nc�WD�i$���&.YR�p�	�1�u�O��4�������7��$X��r�>E�c���4�GO$�KQ�w���4���LO�c#�;Gߦ_���5��Ol�a��nW��XȞQJ�l����*e�f��U(������+�?������l���F��R��s����,�|�2�#���	#�Ç;lDk��0/1}^�'5̒���Pf'Ό$�cR�z�[��ҥ�3�+��5[���'��bK���:袷J���<�%��&�2�����$��d|_q��ڥF����Ks��h��z	�Fl��)ڂg*0\,*EBvTr] #0!�
Q�?o�˒zWM�$p춬�ٍH��#�<�q����NB���D�!�JSOYIW\x�g���ґ��V�:���:w�a1��]���L��O*я@%h�@_lH)���eol[� ��XC$?�C`�[�'?;���1���27�b����5v�ݧ�cBx�d��<�4h$����k��3���<���Fld��_�\ �6�Rυv�6,���rQF��A�A"v�&D�l��DpIG��f��䶍p�VoI���V}�#ǫ0�Ǳ��ω�Ȗ��l
q�?�@dI���(�Ƨ��|ظ�=e�:�)_Q6[��u����,Iv�yܒ?�0���!T[��pz��{��0b9g���Kp:���N�b�x� 9KD����L���S�Q8��)6{���IUR�z��b����f��ƆVN��N}?Ͽ����j�W�}#��.Չ9K*�e~���l(L1�z@`,�xh� }Pӡ�T����E��b�J�~��ρP��<���7���:%��>a��>�i����AG�l�eSv�э�쳫���'�&���~J�,�TΞS��Z�y�%��������beo�Ng��s'|��y�!�t�Vӝg�R�ص'J���{a������wh��J�u���^��X���7��L�JK��9�����?ۼ���Z渻�&j��$���Ͳ$�\�4�VP�*)VAz~7ez�$����f\�tl��+���ڎv