XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?BA)o+�}�,zP/Xf��g"�����pȇJy�b&����п�t7������B>e^Y��!Ͳ<sǧ�@{��_5FJ3����K�l~l�)��$-�nq�k����T��^0���X7��j����hֶ�s�����M�N��m�!���х(*d��1� )6�.uf��{�{��	�7^ɎW�0h�*��j-qͿ�I7�{g��1�[⻬p�LLD�qǪ�m�-r���aU$���ܷ�b,�>�yI�֨z�@��$���{/�+�b�`�K��A"�:t�̣fl������$L���YҴK�G��Dz@���L;v�����z���F_d�!6}x�	�:�_4 ���0��j��o���C�q}_%�\wr��v�a�Հ
.;�\�'���� ��ҋ$(�uH��v�v]�' �r��+Z�ҝeTʶ��Y�|�@!X掰�]eR�Ӷ�$D67a2`��A���`bC�%tI������^i<:O�m6NZ��KlRs��Ҩ�I�y�2�t:��y�"A��Z�H�j�'x>`(9Z��Y5!}YO̴�r�m8���a8� ��3�h8�,}ۜ��Q��c�z���B+�]� �%J�и�������c��ʩ3t��6��s�_��x���5W����<s9A��8xf��/k�$rd��0Ӿ����̄���&�������R�Ex&�!���s�u!1p��ʒ�K��t��Y.3�@]|b#�a��L�*n�I@�Wa�g��4�6?nay�(NXlxVHYEB    6013    1460�"�o�N<��~ k]�N�� ԉ� -N��ץ����8�o�3���_���`��᧶c��u��G � ��aNE��&:L�u�����-�>2�3;u6��ҷw�ş,���d#�	�r1M�����v�ln��i�����49_���^���*�Ť��I+��M�ִi���Ө�h��2p��y:��K��1|�wUTBJN� ���$������� �||�ކ�BN��)�ы@���Jɐ��=JZL)Vk^X\�5f6���MP��z�pv��z'7�G���L(��,��L2�'�;w��H�j��fl�i�y�KV�Lд��9��$Ј�:B	�����>	�@P��D�Z���;�/� c`��Y�)d�|��Y�g���^��1Y�7a���^^��:Y�;��\ݑ�lނH����q�ޓ��>���R`*�sS��m0ʽ�����hP2~�H3E:~�蝃��l8Z`� ��o�pg�N0-b��w@�P��Ki�Q�쀹m�o��G�q������jZ>����@��]-�1UL����^�6-r��w�A��+;RmĹS(�����y��Q�X8CJ�?G��<~ ��ҋ���jO�C�N��0F�J�|e�}5�[:ۖ����?�*�ϟgr��(?&څ%Z�֋�?�OD��('�7]���}�?�I�U8TIܒ�8O�lҜ��y�D�1{�J�x��d����2`��y[���F��1�ޣAҊ�3�{���I.���S�"�*�ŧ�/�8)a�}-�0i�-9B��$m(��Y��ڻ�DI����P鉂�U��_k%=X�J��[��df��U���Dۊ��b��&���Q�����y`�wjp�K4�ւ��D���rdNӨ/� ¿-9�����$�J���#WpN�*E�VD�)�U�mڿc�lڰ�e��ꭙyϭN=ȳ���!��V������]OrJ���Ƶ&��4�����7m���r#�Q�J@�Y-��pFqb`�O�[�׎�O�-�#��"�
U�rVY�R�����I���fS���#���7˜��
�x�5�����f|r�	�o`�&��8kىz����;��1r�s�¿Z��tQ$0wm�@�gt(�U�v�}Zv�?�w3���R�®b���K�M��^����YQH�S[1P\>#.�J�� k*>^4*h��5J���E���"=F�� �հ�={(x\esj�@EbyI��'W�������_��..�)>Ѱ��؂m}��>[Sh��(]E��t�Q7��V$�k�f rAqf$����hX�����;� ��zb�|{C�|(%v����K��y�\�8��[�Eb�q��q4P!a*��^Nu,���O�#���r���߮uA�NTe֐�[���V��U�o"�|��~����W��� ż�����ts�ǫ��iY��͍��NϠjp&�+�-+�2G3�i��k�ю/��R�>`Z�Ȱ������xdi�����3r g��i��G
�x�(^��~��**HiS�GWTH���EVç�?%����>���@����юf�t�1��*��2��F&�ӹ7��}84	W͵/'Ʉ6g�7��	i�s|=��|�7����%&h䞩�����uA8.a�b���cA�t0D�2г�(�	�ء֞��N�Bw���~�Q��q6 /W2Z	�vJ N�p��#<�f��H~!۰)�M�Ҕb�����bg��)_�����8L�M� �&Ǡt@��i����,1�˪z�t�cYS��V�+������[�d[�>Β�
�I;�����0�F	qG�rhd��1�D�
wv:(A���W�>$�I���Ub�cV����s�}���T��+�c�)�E�s�Ԟ������$�"���u"(�#����)ܗn�5���B��8� Bw�O3�}s�d�z@nJT�c��מ`�6)�$��ِa�x�Ҭ�Se��� ��`g��t�l8%+����H�hk�&�I�ǉ4����6�1_�f���ь,	 �傗i�5qԩr,�/���wp�/�M̱#�y>����*�#|b�w�2��w^�ܺƃ�$Q�;sl�����e�0�䓀f�[�z(��:�/�{��05C[�Kj���k�أ���hSWaۚ҄�!�
lJ�X#&,��s�>�S��.��7��!�~���ˁ)ԅ{��Ě
�t���βuj������ł��C�e ������X��E���w[(2��W�-%9:�{�|�)�G6�����jkӝ�Z4?��u!B˺�j�@�=�e��*!!@N�ꈭt]n�aռ�5����q:u��L(����ȩ�cx�@ӫ�jbl�t�!Љ�}]\�Ԇ��-U�tRz�cLR.b6,?�.���Q(/�
���%��Y����^�lϛ_�$u)';KEw�7�D��9n��D���[��ѭ��C
���SW���Q��W��e�W�޷��Y��:BB�hw�����	Aa�T��ϡIC�YG��La�ۀI�t����� ���_�0���#�|B�N.�Ō袃�(�"bo^��m�"<���}YGr�������c!(7o Q�TQ�!C�9�#������؁��Y�I�땵�M�	3hz���޸�yj�{Q����b��Y��]�x��	�X�Ȉ� ���#5\������� :z���9*��[r�
�tG%e��qe7�z�RN`�YN��I?]j~�l��;�4��P���BS����]APH���1-4���
�Y[QA��u4߭bv\vj#ы�4I��W��w�>���6�͟�H�U_,�i��z��p�P͖�D����6Y�jU�]������x�ZI�}�CaTk�[�� ����!4뼄��]���#]|�x`��c 	�vi���mÐEY�.O��4��n��l	���DDy3^�,��컷g#����9��݉'e����#[�?�@�L�Cp{f྄�W�H}$Fbz'Fs��uAh���}��D�M� ��$h7 Te�X.�p�k��UA���&x���0�.Э(���a��]jpY���$��O?�N:b�ٯ?���j��@pǳ��*(��&�f�>T�Ia�3{�T�-{��NV/~N����μ&$�<��zPrI�2�GJQ�qH#=�X.�����M�3�E`��0�?���F��M�P��$x���fճ�|�����#�}�R��HS-�h��ޔ�
�k�x��4�n�c���{H.�::����U�Xɑ] �A���H�Eb����u���	��/'L���ܢP��>��|��9"�Qr�7�����7f<�G����~�r��!���8Xp�d�0���-n�,.�P$a���3p������Mh�ٔEU��f�#Ͽ#H��υة��̿7�^\ĬL��V��jL�1����rz~�s�2��ƍ- ���/x��x|'q��}&�bxN�B#:�+_�U�u�%2�r�}�-,����Bd�g�]�1A�ʨ-a� K�c. �/s�{���cP���2kt<�Ilc��+D	��ƀ�{׺���|��ƹ�L���^���f3���l�j�[-�� �4��t�[� �H�'j|7�����Z�?eT\�'V���qW8���* P���]i7ۋ���=���ohj�`pg�yh�Q�5�#*Y�sq��zEg��Ki����	PZ*6΂���VH7���Wv��g���8�/���P��2�U4*�E��A�CH�x��/nK��~��NqGo�Oe:���~�!mѦ���?�'�Ň��YsS���d�LGo��jf/G 2E�u�-�^�2T���atK�%��ט8�D 14@-�05Kz݀-.u��U'�c��t	\v�Tj���t�k���N!�̥x�~��\�5m�08~�nT?�k�I	��
%R�s1]͟W�
r���;�.�PK��דj��G��e%��i��S;qCO��[Z�I�
ߕ�F�Q���B�����k܎&�SK�rI��������0��Xs�R�
v�Ԇ�#u�r9`�Z���������.���!�NU2��,��2�E�)��AZ��2|�n(�M���_�2��ܓ��x/����xb��$��;�(=�"���LԥR
���XFZ_\�d(�̺MQzd��bZ2�Q���;c~k_��6J��(�6��b3��heSK��d?���"5y�x9��Vk�����/��tp9���n�h5�@}c�
�\զ���:@YH�)Ws�C8>���\C����Y����1n�.�-��_OjT<���/�w)n����uO�$Mr����cgc�|�Ub]��1}�qޣ������L*ka'��JQ�(nc�����A�*���C����v﫰��DI~wk"p�#ݑn��h?~�_L��\6;+����l�LJ�3��z�:�����ݭ	#�i�����	�:]��jA�Dt\��?Xd�n;�=�E=М�ط�?~8�zAl\��F�.E��Zp�|�)�\�j��v���!^("��\�|01l��>�����j�+m�Iʇ�<J��r�01�u�~ ��v{�����( ��kQc0��O�斴�D􄷁���tTt�S�V8�?v
,����hS���e��L��X��pR�:��-0��+���Q�z��\�~_���hF��	\1�Q���G3��Y�}���?Rd��42e�Ї�:�d�Zd�bF��H ��!�����G��CZ�s��*R[k�)�J=��&i"��VZ��������{��@BY&ԑ��kG����'r��2w#�'��#㕓$����<����^��E��n[�nܧ�7���FvZwTlC�*N��E�vHf\3}"�f���c���13�܀�:�i���t	Y@�����5���=Z��u�]�Qt��{>����Yiɭ]}��#�Y`E�T���,S������W��!�U5�y�	�c����U��KPR��[���Y���/�b��hs���<�lI渻G��>&��F8y��gsC��2EKpA{f&��7q(\#�j�ۍ"��{���ŵF�?�C�?9<�R���:R��h�`