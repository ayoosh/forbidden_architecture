XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8�t{��Z�V?ŭ,��┨W�[�����L�#_+����Q��ia�����T������w�����:�_Y�;�¡j�K=k?��`^܋s��:��,^NQ���Q��5��-�SѤ$���O��U޹��0��V�����ё$~�s� �S�UF�C h &���![���f�%!��+c�Kt��?��F�WUm�u���i���ΨA�y\<,u�,T�1p������c۝È�	(o|�����	�@�3�ys�1�ۨ-vϪ㤂o�,mk,�w25z�"�������G�����7'�h��@-\�����6��q�R��myq��ik��?u�	'�D���o�2�}��3+�YԬ}	�LP<�=�p�o"�����ҍ����2v�nc����3��Џ��ʍ��N�u$��$od���/����ϯ*g�"�z��7��r�@t	�6�5��q+�G�ƜV��W���Z�Y�	�˾5�8�ˠtq��e&�XȆ?��H���f������@\��Q�zZ�'��7��J��D<Y`��#*�XkZR��}ڪ���hg�K�w�	{���DOd�,%̏�'	|7��q��h�L�+k�������Q{L�Mviv���7X�������2��yv\`͹�]i�i��(	J��ˡ�~�ˏ]<^��w��7�ͮ#A
1Ip���Tњ9Z���=���i���#��$z 2L:���&_� �dõ�,p"ږG՝s
�� .�YzXlxVHYEB    9efe    1be0�����?'���o���,.�M�{
�	:�^��=ג�6 ��0E�|�����v-]���L=SK�!����� "zx| R:ˉ�1@���6R�!�	�|hU,���N�b>���S�+p��v�>�¥ے��cU�r5Bm]&O|�������U�j.���X��S���'�� (���.�z�)�s�o��d�zt�$�5C��fm>�|KǷϧ¤Bو�!j�3��O�V�����m�d���:k\Б/�շ|w�a<�q�1���S�{)������"~�Y$�ۥ���w2[�G��4��O<G� �����]�mR�k�c��p#K���I/��Qt�����ŘsZ��������?/�ӎ*9?d�2b���?��cJ�~37;�vJק��Z�׿�8�w���7P�:��$>�����6Y]��Q�2t�tē)��u��owÉ:��Aߦ����WC�ۂ%1��q�3|ݞ��2��ܗT��ÿWT��n`q�ᚶ��ntS�]��ѕ���B�_�����û�+8�\7����1y�eYM���o����g~��4 M�e�Ive�����T_A��v�؆@�L�i6��P9Y�*T���K��JY�� k ��~�+��[gW�<�$��wJ]�E�S?��\�����6����/fWQ7�eD��3�Kʌ���Gf}@�[��i�� L�Bc!8����"%��`�ۂw	υ�w��Ѵ��@� �7.��a��J��-:���s
��,����̈́}ɜ?B�b�AZ���(9n�ָ���9N?v�`�j���n��|�oǄ����ҽ��~�X��K��}V@p�{ܗ��yMx��?�2���O`e����9��ZuN������}�g��φ���֊8���u�Tw��{�Z��^�3:������9X�չ��AӐ~>����"�4��O��]�Oڑ�~8�GT:� �5RX�0δw�p�V-���\m��?�}92�X�=����Ӳ���D����vrc�dB5V���OC��	*�g<��0(��u�\J��H���,!2s�uR�/��
� z�Z�ԣ��v?��`�^[�>�;3�Y����v�L���3Nq��~�R�G5e��3��ʹ�jK6%vD�5���z�G?�9��G��������zZ�3v�gd������%����B���A�d���x�����9*���`:Z�h�q���P5��:�my��|ݘޠ�p���e1�0kHᕒ0C,8��$��AӦ����?ٖ?X�z!oY~�T �@H�[���SګM�1��a�LB�_װ04�%]�+6��#ANc���`%P�z�H}R^�/�x9,�JT�
YX]���[	���4L\hd�'ae�E4��!E�}��T��C�5�����M���n��j�?��	����8�]��s��J�W���Gi��߆�f�#�X����G�#���:���FQ���!EIb��?X��/���1X�]7ͨ���Q��*��Y}7���k�|��:��Io�7����8BS�Ǖ�"k��S���9�LM���W�
��%��.��@E��e.}'����ս�蟭��!:W��wg�#�˺�G��L��q�z�w���a}��9�6W�/>I-�L�c��Χ����ś5�/�Dw��c�c{r��ש�1��Yn�������� �p�N/��z��b��n�%KP�t�C�A�dY�����[m��e? �E�Z���N/ĵ͡?���k@�#m%Ó4a�*�.s�Y�Ê�^>(9��WzC���$�W��f�Mv����V,P�en�0ΜO����γ�$�L�{_3�vm}�
L��Pg$^}�[>�L�lJݴ���5�%l�%�LB�1k=�����fY��~(��_�Z�� �a����i���m���Y.P+�?6wӬ��|�k>\�F����O���~����"�y���;=ؤ�$ iݣ��ҏ�(��d�x�B�:���5�'5
V���m]6�	!5qjX�Ck�r :��ƻ(`����	S���ޒH�!Ȍ�i���o7:���Q�m��,4���z��qoПhoh>�3ԗU�*�W{��	>ŉz{�oO� 	]T����q�����ݿK�ε��A��`�ۛ[�P�UNZ�%0�^��&/S��Tb��H��;��/���2���	tOW��7�dھ/�뚧�s�<x�̫�z�$��S�4�XFy-)�g��X���D\��s�`�c�ש΢�?hnNն�`��g:'��}�Ht�}�����h�A;yC�u=|��`��B�i3c�&�\���њ�而x<��!����J���6�Ħ<e�d����<$��I�/l�� /��{��A�&�j�C����Y5������}�_�n��Ӯu-m��^�+��?G�l���ZϩVJk.]Ș/�ة���$��eA���YA�
BF��T�*U��TQ��^x���Z��=U�>���'G�\K�˘�Y�}N+�՗涷��3�3��n&�D�,�� lyk�(�uxa��86��4=�k�
�'	�M�p-S����V�UliM��mN���ϔ�L��[���j&?�JW#Ε�Qa�Bu���X�8X�r�`�bXi2xXAb��C������$ҧ�rU��WW�t�D�<<��(��`�q�6B4���B��8����ó�����u��y��rB�U *n����.j̇�)��ps�i� ߴF�;r���N�$xU�2V�(Z��ۤ}@oPY�`�9�.�J��ϵ�lٶ����6�d(r㒞b�<v�I.����n	���&0;Um��I���>�(ǚ3���4dX��7:��u�'�&�N�gJ^����\04���`�-1>9��Leh��g���q�2�q����}�=)|�$�x��1������/�����E���6f�h�8ڀ��S��")�m�TQ%(�w񁉍��`�5���ſ�a�?pc�K��X�=�b�VD�A�|s�TF�t�9�A�r�q&�us6���I��$�8��l\�i�\m��8B��_�� �!	8��"m\̨917�u�^�Y�C���
_�aM� 	�P�"2��а��9��L�������X<� �SP�>7�7F6��h��`}0Y$T�w%M��K�;�E�`�����-D�/ȍB���Q�>[����a(�]�
��>���D��EElA�+����k��nX%:+�@�������޲�m��$ _�֥�s�Ue�>Ә:@/5į$�QL  "��Q�	�cg�tIV�˰sץ���kK��$��u��X�"8
��$$��}#h���H��K��7  %���x���O�Ar8� ���0T��G�(�Kלᇭ��Z�t�`L.Mw3����[��jX��H���h+�[f�lm4Z��kO&5�n�&]��V+�~чPo�8S�[d�۹�k��N]1��FJe�u� C�Eq��%&���v�MF����E��:��w��F����~��~���H�dB�.�A'�߮'	���>y"�5͚���Rg���F�	��;I+���{b�� ,��~1'���T>)�w2�9����8��ݯ�/�݆)k��Z�fV]a���V�$�Ѕn��F��^�M�>���Aږ�B�i�ʑj�6,}ň�L���y��?./Q��,4Le�HB�%*/J����pf�}�=��f���)ڦ0;ܯY��ţ�Ņ��uMF�CXPm��P�_��\Ջ`&Ƀ�)\��������Q��y"�R��4
:��Q�� 1N%����~V-����D[����=�mχ�=k��
 v�K�׹t�\���굴�8��N���i!����]9�خ�F}�G&�7)xd���]��|���ԗ?�����ͦe)MH��3I1S��]�5��VZ�SMΌʈ�e(6P�*��i^��&��
�S�]B�r�w0���m3��߇=��h��!��B�b]�7b~�i�t��=r	2��5�_km�F�a�L���v ��=x�H��}xՔ��j`~�det�0�ܬ�=)�Y|/��_�؜�`��Dx[mK�u�;�^�"���UB�D/�қ�]�t0}5]zPs{��ޗ�=�P!�#��>��A`�s^+�ɢ�3R$/xNKCK�Es������2T�p��h4��[@@Ä�%�(�\9��|a� B��Y�sxS��OߎC/�1N���{G��A�0�G9��KQ�H�I��3����MC�N�%��VT��L��=�3���Y1j�v�O�*w{��o�3�	��ht���
��* �T�޾ˋ~2!u��;E���ϲ#�bh�ێe�aJ�6$T��Z�dQk��Og-�%N�6>��H��=�݊�L�
��|�?T�
��Éа\A8�5�VZSk�	jIV섭�!h��#��@��q:�^�ͮ�k������#�geb�j�E���7O���IވW[�\�QK_҆���1}u4G?ޡ'~�x$�l��$��$�P��p��X��~q�1�s��I�ayC�Z��ܴ 	�"�P����A�`7I)+��o}zw�'�ԥ��x�N�������s��XI|혆6` J�(�A�EK�����\�`��6?��Cq�W�Qd�����r/۶��;�R���ʴkOʿ8w/Y�[�n�$�����wKË p�����4��'��9��e�t��?�����.c5�)��b�u��5A�D�-��R���x�m �4<ĿYuL_�4�*Z�U��f��Q���e�-����lyˀ��������,߬L�No��#���`��/8�-��շ�u�-nW��i�C�p���Yfl��= ׂ�ms�&*V��t�=L�	6����ʢz���y��hW�E�����%�PŊm?1���2+�U��O/����Z_b��6��%z�mbA��71>lªZ�ѩ&n�ٯVn����{�R���}�q ���ϜΨk��K���v	}\F]�bW9N�\l�F��2�^�������8�0q3��]P�N#S��j��c+� ��욅�MZ��Z�-�{��YPMK0m�\Rz�_��.{���O%׵�����=�ޡ ECLT���Ԟ�*���_�hƛiAy���j��6������\80xa�����jP��Aw��aܼ���}0�9[8w��sf�~P���+����=��&�oZ�Ѿu���b���ڑ�b���>�R�y�A�V�!���t�_�kQ`�I�����(\�@6m�5��v���B���uuM��*��A�6ҹz�h'�j���R��u��i�"C���y��Y��tq!�|̳�c�ۮ��BD��Rq�W����4�2���A~��h����+�i�����iM�u�N��, �^I㔉��=j[ �X3��>!l=�1 ^�� ?�ێ��+�����MP�1P��K�&��6Ԗ�$	2�>z��Rl`xɞS���p	�E�d�N�>s���K[���I�b}	k7��_v!���&'�"R����f-��eK�!4y`k��0];J�Y�7,�Ƅ�r�����w�6h���HjG�cTo��F��{�-��������g�wg�M~�[��[$Q.�K+N����a�~����nb|���ݧ����W|����-n.F#���X��/���/�˸��@>Y�߹��k�Q��^@淞2�ɂ�f��A�*#�Y�;���VA/�M��L�������ϙΣ��bs�&n���?�@���G�Ft�6VR�@��|n�R�;��v&�����w�����Y�\�Dhw��.(��3��?W[�h��O�V�V�F*������fWt[$��~��J�kJ9z�_k�m��3��=d;D���y�A/'����DQ���tK�,�{)K,B�l[Vm?ad��n?��|T���~�������4F����uRY������'͢�1�s<c������協 �����G�p��J �������{����i�$~t����V���]n�+$��b��V�h��n3�Zrٙ���S����������������"V�/Q�qbv��Nc���v���M�,+�]�[�MMf/�&��ԯ���B�)�iW�8�5�UD�'�	p`o�Ӂf��
��+.�KjW��9+�B�������������R��ٳ~b�T|�q��4�qj(y��v���t�ɧ�6V;�E�'{���UhJx�x����/�:��h2'mJ1�R�����M\���9���H�y�ΩQ��WD�J5��g�.GZe�rQ���o%��*L 6kT�&������&B��o�"��֔�4�*��jSf�	N�fK
��ڋ[�5�����<��A���=d@�>��q�csiwp�)�UQ�M�aք|�@R�]��������8t�:�*-�|�'y�O��w�G��z�YT����K�Ey��� ��D�����x\�t�)U�ჵ����0��a����L4N.鶏F8���6gxv�V�6=?(�v�HS��	���Ph���Ѧ�����S���tbDR���!jn�,=�ݝ��j�Z�ܗ]n�'7n�Fͻ Uʼ�艇��7ؒ7/x4d�2�53��q�t��;9:��B��"�: S�ܞ��q�;�\+�����q��q�`r��Ɩc�*�_�5�41C0U�p�t��
���v6nN[�X��A��?�4:�rS����1Y ��x@��1�קr`=O��O��^��5[�n����1Z�c�0�ǁن��������bc�d�ۊ�m��zp��HL�-Yͫ�ͫՋHpYZ��d�
HQ:�ƶ��.�����~���I<]VB���xÌ��T
�
)bKjNT��'�ӽD/K%�"D�%�-!/|�]jY_)� q��5����6Rs��Cwݕ��q�h;��{쬡���Qܟ)�EC�������ʆ�R�c{�n��pm��mU���B��'�U����b抏�b `���"��y�YXl�6��v�3M�HO �E��ߋ��2q�"G