XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8��$G�����4�(�z �~x�����.���9v��<�<L��g�c�˫	ˋ$yᙧ#����7KK��㺤ϧN�;Ѡ2t�σ�����y�F���Z�HQ6��0R���wW�t�M�xBT�{���Z+F��[���c�"Z��KDt��5"��M$��q麒��F;B����9]ʂ���z�R�5���b�ؚfT�8��8�i�0��r^��h��Zy� ���7�]XOOFŝ>Z/�hF���p5W���F������`�~ݼ�(�x6O�q�X�$rJƢ�6S$t�AD�b(E�|�68��P���笲��eNrk%]O,���1�I��[��"�����b����n�[�<�6O��Sr�g�}�MToɥ-f9�;������Ƞ�^(fFk�VgC/��y7�cRr�i|$:�����\9����p��N����K��R���:i��6�M�ך��P��~���*�����|A��B��t�ej	��Dw���z~A���Q�g(�N^�F��=x�dU��C�b�K4�x���ǆ���I��i�B�M�����$]]L�T�l�f���-?�uP7o���c���=1����Օ:�������Q��s��W'��+5�]�gq;ks��t�Vz|�qjSW�V�큂d��ʘȹx�Ȱ6M0�t�?c̛rd7���R�qu� ;B���������_��	�,]TY6�|� .�5�u2�eBݖk�s�Z�m]%I9���7q?�~�wXlxVHYEB    fa00    1f70y#�C��?>[@�߸�n�r��p+�k��$؞n@��.Uj+E`Q}�6����f�tZ���[���*�P���`ncN�R��/�e1�����E�є��e@����hM�g�\k&���̶�M�V�
3�L����D?r4�vL����EpO����2��^�BSH���$w����=O�b^�1	Hs�d�=l�w)��m3�Hv���O�ENKh��~�}����t�)��j9�B���ϖ`���0�@��J�;?�Kp��}��>ݎR_Tl�_�5���bOGC�,���2�ۙ�7�K��!������s<F�и�4a�2�����^��q�dH3?��tV���ئ�g�G��q��퍡�����6�i|wPF/+3{�;~^ݖ�9�~�e:]n�\�_f��*��ғRx����� �M���,�����K� ��=a۵?������j7k<��W���AN�(�H7͗���.�'\N�{M�Q9�﨑��R41-��|���p���Ƹ�6!�� T
�tg������×~�$B�wku#z�&P#��v��Ɨyom0�ɺd��������[<��&j�1��I�����<*V�6�y5a9k��!�=���)~kdY@��A[��v�Hw��.��ޒ1��dC��'sڅ���@:u�*^@u\B ��vU��[�sk\�cM�qҭ�o��D�F�s���s��Q��b©+�Ō/o��Q\�]i襬^��5ԍrƷ�z7��$V�����^s�i�a�=iX��^0���GG�S�4ڣ��P�Mh*����=_��n����d���,Ũ|mi&�	��G�-ɸ���K�X9|VT|O��^{�60=��3>�� �)����0��ExY찳�95��k��-�-@;��^5�(ذ_�,^(?�y��M:Z3�r3+-1wv�z��6G��nΚ]aX�z�@���,Ћ�i�gx�-�,8<n!`�AcAl�+>)qL�9�!�/5-�*ϰ�@������QZx߇�n6ƀ�*r�,�/�(��p�����_�WY��"L�|��T�p�Y��x�H�K6�K�T�{�\ ,8�ݭݡ���tkN��Kce�4�  ��7t!L2�T�/���x+�V$L9B������_���C,�7J��W?�.��T��[í3�Ro��lc��% �Վ"%�����1��N}�G�~=m�f3�f���;ͫpy��%�%6H��� ���,���W�e�j������hnf��N�0��K�.p�k7}I�}E�K&$G���.��#���'@AF�u9d������M2l�Q�77���:�����%	��'�����.}�|�
z8yV:�ז��s��Ծ7/!=d���,�~��n���ph_Ob�)�����3�^
p�39�w܍��c$����������(yM�s�)��ø�e��y��9���+_7WW����W��u�=�������cH�Wx����Z]萊��^&��>�w~>��G�SV̺�fu�s��yr��=&0OF�㏘�Cǔz��f
��|����}��S~�jn!�8���]ę6}�>Iɏ�tm�g�[�H��N-��"��e���2���q��K�8��bȝA*�Q�v�D�MRj%����(��l�L6�3~3yłaϔ���g����@�N���:�A���6m��D������?�h����3�4D����r �R&cv�ڢ4��_��)�+��B���O��o����w�%��5���뢬џ����>k��U���%B��0&� B�BO�������J�'k�P$g��w]�cf��s�Rf�����]�����]��gjBW�[{�?f"�r�(��VP�U�ݒ��%���fje���Ox���0�)��Ƌ0^�_���+������$�C��I�&@�<	p�+��"�Y�|��4��1/�w�J�4�y$*y���Q_�v��C�3<�q�B�hf'�t&�{���ݣ#Ν�'�#���`|�1��y8�W��*��{A *V�P�o��ax�;�|����zki����q��9�hO��PJI%��
�@,÷��6��ڥ�9O%	Ε��`��~j�C�unB��:֡���6$jfɵ����p��/���H���&���I���黅��P0}��K:���r�s����b�H��~c����1#(���h~�[�)�K�;�pyx���a���Q�S	'���i����ݶ��Qa���������쉅��	����8c�-��E��_"m�2�O����Q�����%b���p���D-(���<�.�_�]"H��i���Z��4r��Yt���o�� ���[]��SuxV��׉��������l�k��<9��N���u�v��j-���r����b��#f_EU�{�5��C<J }_kEeEF?\yT��t&�'P�߹ɨY ˼���*j�8��JdJ�y-[,�\�ƭ6X�%j�:��+~��d�e������	�p�7[ZM o���A6l��*��D3w��mvԅ�l7��l6w��ĉ��$3��������wʱ1i��_sIC�[�
�	=�������xO0?�~���Mo�޸(w�~/&�L]�y�j��v���t��%����>U�j�;������f/�j�U�.�� ����=�i[T,�FP�<h���T�ԎܹZ����6��:]�_����6p0�l�65[��� ��cX�dQ q��s��Xh���;e}w��&�4/��߆�8z}o	�����������I�M�	�x���e�0���I��kd��6�,�� v�ᙇ�=�t�N~��G&+߲��^_�	��ӯ��e� Tz7����Z0��g����T��ܚ'N��4�z�t�{�o:sΪ��0o���zK�^����m',�
#F����bѸkE�Eg���o�:M�e��0݆����s�z�ʖؗ��� ���;�S1�yɯ���8c�|���Vr�b7��m�Q}N�!�<�!�Ia���&��^n���	٤8�
ၬ��^��\�{;>.����RD��&L�\O�
e+��N|�6�N_Yz��&��.+p��c%�r�Ā�`ٯ����9!����q�����5�>��K�U̿@?p��+=�,�.�k�)��`�0�Z���G���U_եg�ު���Eb�}�pn}o�P¸*6�k��j�ב5����I�T���A��md<��~���B�E?RV�{[a(Gz��XN#��@�M��0{�	���-S."&}a.S0���+��Ӡ��t���<��=��tb�Ψs��~��l�v_l�h}g?9l4o���3'�|��c��%](��vAuC��"�Z�%���=0�N��&�{��`�s��
G��6M���\�02�Of��%�\ǂ|V6QKj�TP�*5�9�Fl���O'q���Ug9��~��\ѱk�|�'���E퇺%�`أ�-��T6n�"~��;Z3�Y��D��ˁ-��@+#����ǹU��:� S���ѽ0�>0���"���4�L`h�L��\\	_����C8ª��rc��1'���p\��o��s�|N���-o�X'�L�z����T׹) n2�' j���"=U�j���d���OC�i��DDt-���<^V����g�i�p½������%�p�^����q�h�Y�2�s�ݝ[�1G��A;��PJ�B&'�.Y�������ɨ	ڦK؏1�m�� �Z��+Ԙ�A%k�/����`�}­�1��Z��'N(K���8oUM�E���4����풩��0,��HBPF����)=뚃r_�À+.*�,�7�UD�[^֕e�q�A���� *;iϖ��V�H�X;=�K�|�\������M�z�\P�5�`�1�/���]@���νMh9ntF�����/�h�i�+��o�����]k�Tސ*U��ё<���(��R���SQD�p��m��>|��ׁ�īF�5�E�|,��]�u0�,I!=�������cl%1����ߠ"���a` Ԇ�9����$�"f��h1���N3�`�33����a�S"^Ǳ�����Բ?1����	��B4���t�yyY�#@=�E�s`7��j+��;ݭ2�d8L9��@��H�r��[����q�c�û30SS��ت��w!�����F����Yi�o�c���m�$��=kp܋	�4�6���1�ٲF�	�u/8ظ#s��J� P'?���!\��F�Y��d\;K���q�wu(��*��x�S)�{�Ҏ=S������7�kj,a7粧���W�hH���������h�r�o�3�&[�M�$3���t������>��ʃZH���8whd�K߻�c����tɎ�݃n	HzH�uT6��\���M�MN8�<06���!�q��/�_�}����n�[�t�RSY#
��4P>v��a���l���n�(J:��AW��( ���óYu��i�!�{]�=P�v��[E}���kA/�z��D�.���!w�t���p�dyg�~��oz^���C�Q�Dq�C�a򩅦O��ESO��ҵ֭�hF��L������C�؉��M�O��˘��Ʊ��*K��Y��;�9I����.6�X�%�cU�̓�K�b�A���H�%�{/!�Y$̺�^�j2
��k<;�T'��bi^R6�S��~��6`�ɫ�m��k�]�ɰ'�ɠ��#4(�	@G�s�(��B/ͱ�;��f�	k���S)� ���:R�՘���e��_�WҨ�����f	i�{�2w�h�_�6d�_��ouh���Wq�w����δ��dv����y���!����M#Yl`e4�ruo�eK�6�	FR��O�Z-���9�P�ަg��JG�rB(���H
��B�0�y��F�=wc�����V���	�T̈́��Y�ҳ/����4i���t�Jy^��f8/p�pV:�+]lJH�3hΤmF�[�X���4ޟ�~*�&
�|�ڄi;Ry6�m(���6�Z���@�癫��?��Ѐ�χ��!�]����0�)�u�L;�MZć��B�T<��u"�p��Q�����_/z�}�0����;ܡ�$7g�GG}V�ҩ�*R:LcorE�1Cr�.P���a���̾��46ץ��	����g�]lM*z�7��R���V/��;�]3z�Ԑ�;� �W�z�K��t����T��h���pcݎQ��d�L{���@�/C�[�bE���Q
�9�ײ��\���W��0�%�1Nq�<��#������2c���[�cj�X�z�?�c1�\zǇv?�Z�s����@�E��!͐{�<�>Z�d4e� ��Q���%��Ϊ�5����������7 b��	��+�g@d��j7�-WS�J�2L��ő(#sc�R���"yz��b/���o�2�p{1Eu�6k�|�Z<H��Qюk��:Ѡ;7WVˋQ<�r�Ѱu�E��IH���]�v1��	Cfy��A��a~��p�WRQ��Ur���J�5�ke����;�|O�څ��0�aDj]һQ�X;4�] ��zҎ��G��R��9.{A�z`�����#L�s I�A�^��
���]嬗� fw�}�U�X7=xQm���[[��[��I~�~�`S��
$s.o�V����y\�cc����������z+x-�i'��*`M����3���xd}���(������D���ei���,YտKݓ�%�X��B�>����kn��E��-�͹e��m������U*ljv'��?O�-�Ub��r�Ga#ꏒά�I�o|����ڀi�I:	i	wIWT;�N�B���ۊ!x���w�Z�>5׷M\Vp���Ԉ�I�vRL�{�Y)��,���&��8
e�]���Va���pX���q�mg�O�� �܃v��AC��7	��q�"����j��}Vz#��+&j��o�^��(�ޓ��Gqn8��ؿ4i�\�����y̵��=WS+��C�l��S��-�I���}�K�K�')q[�4Y��h)M4XDQX��4�dF$Q����o�G�����,�o�=e3�1<���G�b��ǭ�4�@ﭭd��%HP}�t��� <*_��P>#���W����`� D���Y��Uc�h>?K>Ddd��v�&u���<Ԃj.L�}�0T�sY��Y��B�2�n5��&-�ڮ`�D=(p�s�8�`"�[@��[:iL��վ����`�nw~���c+���F�?�����_�씩�x\y���~v����$�UZ��2���Ϋh\!d�//�7�E�X�]B�hZ������h�\����4uq������O}#�q&��q�����¯Rd� A�Yg�\Zú�'�*S���N8-�u�����IKf?���1�b�"��Y�_~?c�g�,���2��
�}��gr�l�T�fѪ]��ެS<�7"�B�ޔ(�g��vR��K��w����VX�\YOU�G�x��-d]�&Wڃt;C0K���e��X�β*֢��@C�v�'���A�W��S0iA ��6�ۿy5h._�=�㉦�{Q��b�[)����]03v�]��y�L]�Q7�a�<��?mZ��� ��'2�'�A��{.e�͡��K�C#��,Q:��>��'���6�W�WO�=��c�sB�{K5][���챋4ed*�@��.�yFäY'S	N�J���by�ʂT�N���8;z�����ka���&kpc�2ޓ;���`�:���n�%�gK�})��dú��ٯ��c`��]��!��|z^�����!.߮!�Hu�$��t���ę�~�b^�|���H|�z����օn�w��f�gӱs��������i=N��<R�w���W_���o��V������J4�n7�N�:�uA�ZEP�D�:�Sb2�����V.����R���e�k����FVs��q��re Ȱ����aD6B5w۠�.1*��YT:�2�2��Wa�}�1�^S�P^��\���G��qH��rw�
�.=��G��vO*�l��n W��C�y����GR �2^*��&s7�c���C���Ӌ�ǐ��L!��K�7Ӱ��c�;�ȋZ2�64SD�p��]�ۥh�Ta��׆"�A n<F���f=�Yn �uU>m��t��0�j��/eC��S֘���"�Ĉ%B��}|3
��O5�q%��a9Y��pK����k�V���z�H6�!-\(��+v�x��B�W�AfS�C3��J�+:y�,5�[�l�\�xj�4�х)C՚��·���pCE�ԍ����P��	�+j�,& ��@�CT�Od�;�_r��>C~fs�u:Lz�^�ՇX��nǑ�L������{7����g�(=kAS"��2͛������w���OV��1bI}9)Cܰ�1I�C�Z�ظܹ���Vԕ��0�ɳ� _�u�D�9�0jD��`(�%�\|'�|��K�ϐF�Z(K^;����(��UY*�F�ӒtJa'�F����or��~��ʝ�6m$h��J��Edo~�����6��V�lq��*Q��nj��Ӟd5�9 %��dW ��DA
��#.�]H�Z�e�W!�1U
,wƀ��@A��)<3�i	?@�4J�ﭑT��pe�83�Vͦ�3���pH+�X����v��X���䜆n��K_�Y�S_7��T�o�F$̰��H2��~N�֒��p�h�(g�'�0��/�|��RG�
�[� Z� �cJ��5Y'R#�iu5�Ж+2f�b�IH̹�Z�ZM��v^F�(������z��*���}d�x�-r\�ݐ�om�����g(%i�a�m��y?�/BD�2s�������������?Y�H���W0ݠIvС3Ʌ���XlxVHYEB    fa00    10c0/�������Q��u+� ���=�h���X�@�i&S´�?kU�dH@E,&kke|S���be��&=횳.!�SO'U¬�s�kwe�qt�q��}�#E��qF@��M�q_�X���}�{62еn�mͤ#�d��N�oI�qcBK�2KB��zH�bv'�����&�]�S�Ft��mo�$*4��Xӝfyn��)�g��TJ�0��4rři+�5$����y]c����]�=��
C�������]�`?�Nha@t�F+m� �\�fa߆Ul��@L_)��|ۮ,+���1���\vL��]�\]�
Am9o��+�LT�m�D��g>�Ja�|k��`V���\E��%k52{����������W�YcT8 �/�
�!l�Fyv��q���$t�v�o▕������:���J��mF�Y����
Kܜ{x�N�:g4�\�����]�a�pB@V`xV��5�V���s�W�s�}M�ڱ�?�����uʆ���ƒ��@���'S]�P�}�Z�0�t\�r��e�Z��DG�h���F(����z��V�K�Y�/���c�L% �b��7Ԍ"��	>�)iD�m)�'��D�ķ�g�8}��?,����MPm�*�����Y���ʊx���������Hb��tZ���oC�sp�G��M���}'��s��ov���FyL.�4�D7d�P�Wu���+�7�R�7���1�����dW�.����5-��}��E_GGc.�N3�{���� T^Jɿ�L���d��}.��,l��=���a�	��Tf���d���,HtQ��_ә��;T-�%��>Zuů;�#��*�~ox{-���N���Ɂ�^^�a�tf���ְ�.wC�р�?L����,'*�d�!.��ܵ�}i<��w�f#4��߇>�+΋ׂT�M:N���d�B��Z	�&�b�>�3*6�]p�G�@j	��9G�v��=wūz�$����Ɲ��@G%�(�^5V�r8XB��D9J��9��R����t�ǃ_���"����ב��j��A0t0��̊�w! |�\���\�T�Dq��U�w�5����C��D�WbJ�z��/
�j�D��GrMnq^��*�#�Ⱦ����y��*�rj��A'
f1<���)��CZ���X5*��fCu,E�ѝ!�MW��$�������ϙ^#:�ua�Y0�ʟ��n�@�W�ȼClY.��?��&��v�$x1��Z�I�^1%��v����|^�b�4�	�2q�9g�,�Fč��#��e�b@������@�g��=	���L�ug�u
��m�=���&�<?���0�g�<�U�I�=�<e��� uH1WH�`K@���
�qq�Gl׃h�H'u���x�c��&K1����p^P�H��c���F���w�^�J��V��m�F>cc���l�+q����a4�oc�um��͕����Bd>kW:���Vo���{���
\9��H�j�7,����f�9Y(�����d�c+�����*q>��}r&�j������� .
j��0:vKI����[��`T�.��0powpI^@��L��R
�[b>ш�X���ͪ���֡e����쾗�2g�Ch���P��%�c��J������1�����+Y
.�T��ޗ��t9�i���i.���y�!� P�(���B�N�0#9�:���px6&Нߐ8N/q�J�л��Y	����_jHJ������b���U����(!TMЄ�1d��8�w��o/���b:����CO#�U�����e�郉�HI,��f���7����%Ʒ�8�+H=�]0H׏L���pO���� �����,
�|HЩ3�[JP2\	\���O��G곩�g�i<g˺��5��R�:�M�0uN�Q�bC��o��"H;�]��n�%Fk�,"]'�mBn�$����F��~֮
7�`?��L7�rT�5�<R�2�V%�K���;�����x��<���wF�=K"�FUUv�~Z���_��|�x��D�������e[b~ݫKh��N�8L��x�z�+�fj�v�eB��S4W�lFoy�� �0���!�[��H�q���f�m���4�B�/���P>[6*�1[�1�v>VQ�d�
�\3�_�V�٢��p9^%��2n�4~���x;���M����_s��S}�]�����m+�s.�!j��]����l�D^y���X(��U���RP�d�2t��4eR�V���	�ۯ�W�J��e�M�ǵa�?@\�:�&��Qm��Ʉ3R����>fB�X���8Mj��Rd
�Gc�v���)ճ�:fsr�����"U�2���Qܚ�	-��_�l��2�X؄&� �m�}�Ty��f���
���h��i߷s�a!vt�%N����VP���!��9)~�+o��;���Jgޢ��Oem���6��|��	[����^ڊꌨ�����+4p=��'��y3��H
�s��Q���E(��ѕUҞE��.@M�������xUKe���G?y<i�ŭ���2�5����WH��?������"�����~�-YDV	P��K�6�i�ל��� ,$��fιqu�pw�,@J�uC������S��{��^SPj��� .ǣ�.�i]����Et�'��ɓ�e��=?k�X��0�9`���/��;��E�}���tSQ�o��U�`	�����\���+俧�,�B�{�%u������Iz�l�����~�)��,E��?jk�X��:Lp5@_����_5�ٱ�g|$�t/������C�%	"�?覢%�jӞ�'��wC�/�V�/SfXB:�C�iW��Nri�h�Q��;�����C����>�[�\���K��v�º�_��#ɶ ��I�署�9V���d	V�<t}�ҼpPw>�+�~L4-����)ЭEjC�`���xH{e�ܱRp�%��+p1�FN��]�+���&i�^�I���7|���Q�I�<��U4��l����t���r��4\4��^;��?6x��,e�5��T�����f'V&$��ߖ#���	�+<zV���Ɣ�����H[}�D����n�j=�����Uy��mR���>ߓ���_F�-(�;��D��4�m���|b������|>�/l{	�!�
T�,��-7D۔����F�Fu�z��L�n���ig�!i�M�5ڇ����W�\�2x�M����)j@1�u~��'���>��v�(�"�q�9Ævn��`�B�!K���b_��1�"��'In�]���� @�7I�'�9V̰���ʕ��9��)�4��%��Ĝ~���EٯA�o�Xa�g�f��4,�f�� �-'_����SFEz,/�1�SK'���U�Y�`�a����-&���>�b�x�{U�B�]�f;#BI�sz��G��94���=�7Q¤i�p�J�hT����\o�/�.Ӏ�%p���)��xG����8 I�V�,4���Շ�x�AYʅpFʷ`���|7FG��V��I&Y*�r@\/�4;��8^��ݐ�^�a�6D;�o�D��Ϗ��jt�)�\Ml,�2�i��B9@����%i#�c�OqC4�|�]Ll�SX0��^6�X���q�ߙ�a�&CmI���W��2�������|��_��=n�mT2Z��;����뜺n3�Mdd�
N�M�t?ܤxO_W�����вt~c����A<~�����%kqa�6�b�g.P�fX����<��0�ޞ$sr���h�����a���=`�5zO��,��`�cp�����q���>g�,+����5��ڦ� _��3�Y߄ޥ"�}eoY��GS.a�4�.����I>�)�nX�����B�29{���-D�3����=t�_2�����m`$�V�{��D"�di��(�nDn���/$_�t�vݳE}��+U��Zbi̋� �����[��g�n�'�Ӆ=�l��Y����J:�D	 o�6�op�j��3@�ߢ�,�4u���-(��0�X�눺�n
F��'8\�{�rr�	G�'��6�=U3���ꆸ��h�:@(�f�*͋B���qtE�`_C��s<���Y�d���%]��)l;�'��iM�vt[�N\��b��y��[U��]ͺ,VX�w���h\D����i!�'��U����0�y����_3� �<P�?��^A��Jnz�]���\n�C땰�XlxVHYEB    fa00    1140Wcr�9�iʹOӟ��C�D�_A�ۍ�>8(��7^F���ӷ��4=$��̭\:Z��]j�9�]�[�4���??0^`�}�����n�S�r��0^L�O~�z-~!���� N���S����[J�]T�L�|N��	�Zwc�?�s�� ��nN�"�Z'T�3���ё�� !�� 5ZL+�pe�u��'R7�����	ʴ���e�:������F�%A��ۨ�}�b�9���a���K0��ӫ��?d'��w�7��.bWt��;�7ӕBSS�Z-��c��\<,����}�=�0N�h�2o�A~f
�����BD�Y[r/�&r(�y/}�`Nu ���_�b�G����;)�Ghp��_�v
�K�����F)�s@ͯ��ơ���0/xD�J#��}�t�A�����߳�K��Щib�
Y`Da�o�x��Jr��� ژWVDQk_�������Ժ,�;BCL����	��A�:�ѧW%%'��R���7�� �����N���Kb���W6\ P������<�����������n�|����Gѱ�6v�/>�(�^����Fd:��ܻ_��(�X�~���Jྏ��&�>���[����hJ7���y�<�3I]!˯P�e�9 r�)2�������(�M�fa�����Њ�]��!)���X�Ou���]�\O�-���&�i�?^�A�Ų��3�[�E�4��Nwo��6�ǟ��6�љ&��N�M�҉�@�OP?�aWaq�oY@  � ��UO�,O� ��7�s�Dc��/(�<m��E��9�e�K��2I8���nX�^�>�ږكBP/Ib4'2��~K=�fL���ɱ;�P<w+d�	!{�k Ǡn��ь"Ev���b��,t�Qe���75���=�/�Tx�!��
�y��P;�:`o'76gu���i�����K'K�ω�=��!x��]��a��Ҵ�I�stq=��!L�pt��I�� �~���T�"�4��]�i��gG8���j�[�[����@��>��66��(]��b*�u�T�&��E��}�:�+�S�C�Vf}O���v_Qw3#-�{m���hH���o�Z#�P��!P%�㭎�/�2�����ܔX���;�mĬ��~�놞��T1�à�_�eo�q���X��A�\��Gyx���ɶAF�{j�'�:~b@�8H#�ti��M�y�gJ�V��B|�Ry�6<K�/+��1�7�p�w��">�ՃӉ���,���*��9Z	����cI�:v�^����^�O=9o���21=2c���o�|2�᳘]�� ���#�#�����^%�t~��7���`	�>�X+ �Y�����*�[�P��l���Fp�k0t�˫��Ҙrg�j$ ���o��6����_�ʌWgw���VH!��d����`�Zh{vLT��9�N2��⹐�{��M�{3��(]a��*�96+u�!��?�EdC2���H�K,lVGn����ܷGD�k�E��Ug��&N����?a =�C�/\W��3J�㐌DB��#���K	�b��.��?l�z���֑{f����vn�����׶
��FW���kΘP������p������z��?>M(�����P��w��[Wd��A&ܞaч�Y�I�ԥo^�ʱĵ�� �ބ���$v5���ᚂLbi�%D�δ(�۶S��c�-*5��7�+("ܸ���9������]�$��-�&)Η�0��!�v=a_�� ��7.}���u���q���6d��Ĥz���ul0�Ѕ�u�0gs�4��Uv9�Z��2�H�'p.$k�K�I�����$�����bu� �fC����:9�`
g�C�%��4����e���?Ol��M�u�臰
J�{�Tљ�u�P�6��&�C~��ʘ��F���� ��avJT�<�j�r褕N�	��SIs�ڊ�-�ͻ�/�o�O�K��3��c`*�0P8�%�()2����%
ssR�f_"�s䨩���7���ZT�9�q�Qx�qC
�U�B?���X���|8���1��U�`i53���V4��{�M ���B�'C����'[�C�pY��������XQbvD@+G��w��6������-�\Dl���7�&u��e���>4BD`��g��m���(WN6�������,�N���s�d;�>�8�e�}ew
_�9�4��H<j��ڝ[0��9�:��}�p���\����`9-��z��bF\'�/ -r�,�L�z��"(+��v��]�?���ې���!�3�7�m��$�4���B��6�T�	�#���1�scls��sG6֜�C�r��Ù��?��=x ���Z�Z%A[����Dͪ=v�*Ư(����e���̥G_!�<3�v���b��a�P^�#o�K*��W(E�'��e�r▷��!`�Wz�
���yM��.so�r����ڲ�_G��A�3��}:�5�6>x�0���4|���_�e5��^AɁ9��C)�A�GUZX#�q���D�L!��J4�/,<"a�\��.;�GY�SB��(�b��he�E%��sM���n�����Z��-&���� �V'�9Q�j��0��ZV���T�?�'��D�4-�=z��'���nN����ݗB�+J���;�����8bu���v~4��MC�9�6����D����28f�1a<�x>�p�d�Z.R9B��k��4����Pw�4��Z�gEޭ���x�n��+�Mb�bDnǻ,��e������P��=l���~U���~��[����E[�K)nF�L�T.d��<�J µ�3�K�/ZF���X���Ⱦ��ro*u�S7��� ؄����7�b�ԮU--hdt}��55Qg�͏�V�u�:� R�s�?׸g&���ޮ�PC����k�NB�i$����W��� },��zF���L`��Jֿbk0���,�Uem�}�[�����w��:��*9?V�E��Z���ݣ�bb-���~Fa ���q���rd�'���~xkU]r&
*z��m�96")Gjs̹�"X=\_��!+)�!ļ�i��wW �[G�R�o\GB�.NO�	BRw�ц��5"�j�AB��&Sn���ްC�}��4�-��GY2@6�X\a�|�ZbKL.��"~���2��:f�2k�r�u��/>��2~�	��3�t�,��7Xkt���S؏�*�8j0�E���V&T�.<��,�3Yܤ��&�2Y�v\1�����A΄{E�:������-���·%��1� ��KuB����[�8r(��sH�>�Ԋv8F�iȦ��
��� �n��e�:�qQs{��o5�V�r|,�PC���?^'u����:�si$f���	%�K5��X�B*���4Na9��څ��4��5�܃eN��Lk�i�*�:�%���m���u$��$`��c�hp���N��i�����R�Kl�ă�����p��^3z��__S���KG�~-%�V��;�?.�djT����e�(	^d�pe�M��$�h^��*WUa��O�צcK9]�T��-���'�������!a��_Sk��K��r�����5���aNa��9��H'߹�c\R*'���+/@�wgQ�$\���2��Y��Mq=�jEAs� c�O�2+��u�+6���>i���́��8Z_�f�������'��n&��R�-�1׊ �]B|לn*�`\��|���  ,)O���m��i_L���8�n��-9�}G��b�\��Y� �iB�۸4mǞ��w�Mٜ�3=�D71 ��*"�!���z����KZ5���?=����HSy!R$��Y�_F<�[�+�+�L��ܼ`A��:ǹfv��'b �g�σ22Y�<*����7��qxg%�qE�^H�Z�>b}1Z�����<I��Eɏ�f}��ΫER�p_��Ц��o޾E�A%ƴ���t;2B��� �[�/pj��pUu�C�n&r�%Bb�����_�e�}#����+�}����y��E���#��sٿgȵ��J�ќb���k�N�!�ۗ���[���g�ާk��I������!I>]U�e,�=d�ɉ��
dZ�WSc:��"�f):~���D#��������]�5���+�j#Y�G��y�B��g"�(X��|g42Vs�y�6#p�T}�Ѵ#*����hs���z�6��G܂��6�ҕN�H��*���CL����U�����E�M�|�g��9.<�ۑ�(���r�#����	�����������hCr�O�|������`2T�_4Ϗ���7�f؂�~�0��XlxVHYEB    fa00    12e05Ά�iˀ�H{ �
������i_'��9X�&:����R�t��שL�ly�E�Ţ<_Xkg�����< v?G^)���o�%�?�'~��l�#m��=������Q��>�v�p�W����`�8!��9����xP3�*�;���WyG[�Z��۽�������SE��]Kq����(���$=r��������Ί˺�^X���a@]��w6a�����i��Kݑ��	t�SwX�"#�Bi|���:@�SG� ��E�Ob��P��R�Kr�%m�vz�U��CF�g9ft�Sz�v��2���:���]��S3>9��*o1Nm��j�.
��M)���qB�IϷqg��}����R�(�x��^��;�ab�OaIW�~��1e]��`���L�s=k��SP'���n���h�h�cG����d��G'����J{w��� �K�
�R�XbV�����3���P'� T�Lk�8h�&G�t����Ə�
���M��`�-��y�R�- S��9]�5�23E �����X�=�	@����g�li�C�����lS�JB�8��p��
���7SE%��[������c�rb�+�OR�����A��gM�?  �sf�w��~�PxHˁ��|
bc֫�.>����|	��P��ot�+�i����!��C��VO�">��-�)���P�L��7/y��u��א9F�<,3�{�JYjH��
B��f���6��dt�'k�`�ⲿ�+y	��#1(�o��`���8\YU�>@rk���?�kb�s����#��1�e~e����A����p{�N�2�M]�pD{�ЇO�!�Y�PCZV���}�t�aH���9�~�����ީ1�OTQX�#F�#h�'�%��s�O��\�nQ/��-���}G|=�",�'����`�Z|g�"VÞd�ъ���}���OfQr�KH: ��¯� ��^;a2
SN�8-�0��A>��O�=Q) ��{�#��]ՐS��Rz*����|~�5HFl��\y�W�Z~�X��q����E	��ƹ&��cdp�KVƠQr�\�+�{s%��
䒬V� I�t0s�J,Y�8��yP:ґG�|����[�׮��+T�cN��/���M�'Ծ�8Z���à�/r�K(��U�dJ!�K�]��R�BE��%���U[���%�h5��P$JE�W{���^��>��X��J�Ղ��^7h���~�]u��6�=b
\Vm��AZ�e_���?�Q��Z�i/ى�es�h$�;m��(Fm��vQ�6z�-�r����}G9�}���~e�Z�gWĠ�فË��F&�+�
��_���6%��`s'��%}�Fj�$&�@V_��H�U��(r��G��g������ �K��5��ّ���c&k.(^�Psp�F��I��t����'�#ov�c;ļ�cf3�[��jS���mb�-^���U|��#�/�e��سfX�ݙï}�����V�awa�GaEg+s�pA��A{����I1����dy�Z�QG�v�p�sF����+w2#l��iQ�9�����;U"/�+��T5��1^Q��H4t����#��F]���1:�g��˽�!��Z����ؔ$[���&Ý^0*� �]��(��4.D㧐,-�Nmcs��ق����8�*�����A1sH`��w��	-in:d�:��߂���O⃯��mǟ�,�3�ъ�y�`v�<:�ߗe�|OiW*q4�[D�G�Wb}���쮈\L5�Z�;x��_������R`9���W��;'sB��g����[bQ��o#�|:���BM���L��ˡ0�Z��X�5�~������G~����t�E��:+�3ǽ^�X�����7f�̹�'N�B�a��$�0v���^���\�Y���z(9�?�Dxi6qv1]�D
Ɇ+ڗe�+�:�@?�	�z�b0L�ڎ���B��G��/��:1��f���+63�5�ԡZ���(k[�E�{����(��G��͝k���<�A��E��M������Tg�{����>���E.y���g~��I���t9�i��R�}�49��>:�h���q�����p��n������t�1�=A��} !�O�����X�KX_�a�.�]?DÎ�@F0�b��Ё��z�B �/�d\���3t���m�z`��#v��,�f��v\,ˬq�h�i�,t�P'�
�Dz\�@���Z����Y������q!e��<�S��|}���s���*�m\��FK��r�4.��,5H`:¥Q��Z1��Yk)����U'��$f1/6L�]9���4g��,N��9I-�l��JLH�e����/B��׏��"�S}�C����1���e�d�e�����\�����f�$�� ��̱E�q�s��z��3��"�J�MB���İc��1�X�5�s�DB4r!X�n��u������L��[��0+W��� 9~��ߦ�K�٪Ɉ��������E�fZ��VȠ,�IT7�WM<�`^�/�:�B����+��\D����H�9"�����%�� {�b��ϧ�GO���}��~����FͶ�V����c��r����+_����"�Cz�e���Q�PBF3���2�t��n�KJ]�&�1i���n�#�+���͗��*����aM�=:2�5x�β�&C�u�^���V��"I�n�~�c+Ua�ar�|���k/2���O��C���#Ȱ6[��d�w�����%���ӳ8��v�{���}~e��y��#Ҍ�eq-��kթx �o� 
J������Nw�[ʣ��74�|�Po�${C'� ;�_�����
y�a ^�_�k1͚��)7@]$�f��X g��,,�	�U����T��Gs��Z�ŝ䇱�b�^@�t�&M�k�!"��Hä3R����e���ڙ��̸�2�����'�
�Ǭ���>�ldKBƳ���hO��J�.�@a� }%���4Y�Dźf֐}Z�}ǐf�p3Bt�M8 ��15�������*�~�X���o��}��nA��2 cp+B�Q�hƏۃr�p/&g�Z������+鱥�¬*�{_uK��(�@yrg0�'�q��͠H[����Y��/���!дT�9_:��lp}2��R��gG,dm����Fʜr�tsdY��uQ�vD.u�z5(r�v<�+X�����P��֜<����ɗ��s,$T��B3�x�~@��mL���&���ܪ�i�[>�WB��W���u������_$�Źۋ��Ϟ��N�^l@��ln��銍�{�]#?X�t����ϔ���䜷+C���v���,�2!����䳃ң�����q��3��[����P��4P����0�-��A�eR<X�i����C�)���71M��rB��w���b+�cMv��7�`��@�����(	'۸_�QC(�
G�5��	��#�b�l4�J��t	/3���4h"���><�Qt�Z��Į�R(t9,��B�-��������M��T��ԅ�.֚|m�K8v�}���Q�O����u�۷(���������iz؄�ǩ.M�`xqT�^?�C.[�Iy�G�m���G��.��D#���0��D,|�S�؊�h��V�%�~�J�v����Ya��K���ʋ�Ę���}�h��&]���Y +��ր�q�ܖv�ߨ5��#1��=�{��ߟ��K�,Tjso�c,+4��>:t�B�=�!�j>��o�/����R%�˶�����Aa��Ws�����$Q
.�g4���R�����j,���;iV�d�[��!��0iP{ٵ�,o��!�H��S�]	�_Y��1�c���ޑ�u�G�|ᙱJ��?؇V�?O�&'��6��z�*����������
=n��T�t;F���e�D�iц@M�dڅ���1#���~xæE�%��0���5�>6��y g<��Tr�D���A~C=�������g��F�,�#[=���0ݱ� �x� �7K��n�uJp�صC%����������Χ'J�.��`7���=�������[t�A�r�������Xh�u����ւ i�0I-����D�҂�zU~0���i�+��ϗM��������:l��[|�߀<��+&O^Z�W��
@w6%)S[��e$1LlÃ`� �T���0_b�"rD��ݻ�u�W����^�⿙���<�,��w	8a?��\o���j��a�d�)b�-50�d���P}�佗�+wXW�U���9 �D��\1���2���+��p�V�4�zx����"Xq�ߙ�_�l˦,ї�ݗ(�������B\��/��C�4ć�l��hg�CRI����ZQ<���@�q��,��vy��Q|y��j����0��̋�H�C}� ��"�JON,vl��)��&�M�7^��i�K;-�2�#�<9$r�>��6��p������W�d�K�TeE]W|>p	�o�m�W��,�t	U����	f�
���>a�L�������" �i��4�Q@��Sn�{kfJ+XP��r͉06+/�H��k�>�N0����M6	V36~��Hj�.��eFGf���~���'���ʨ(�7��°u�B%���vrݚtR��Il�0}��Z$����[����ȡ�T�d���~_�+�Ds�����U �O��߁��d�3�e�S�(^t���?�#�M>�g_�-�~Gs�oa}wpXlxVHYEB    fa00     f50������я%�։��O 	�>�Z�dP�Tuo�l�($!\J.1�����N��X-��9�VV˃l{?:� ��#jQq)���׷-�?��ꨳ�4�솁�j�l>g��Z(��4��лFq�y,s�!�Gڬ:!�U(�t��%��ru9�R�~4��<0��/ �@(��_�%;��i�f�O���=E�S�7&WTI
x|'��
�6�-?ﴇq�oĠ=��Wi���<xp�<�ӽ	u�bJ�X[mȱX�2��8r�b�>6E�܇�^/��\�0��@�:�
���]J���?*��Rt�C+�2�b?	0Ⳋ���y�Dj0KBZ�Z�K���6��=����w_)^l�Ć�p`��Z\~]���`�������p��p���6������vE��Sv�J�����EdХ^��DGԵ��XA�3K�w�ΨP+��B��)->��0#�G|�6g��˓���	� �r��&ν���!��K����_����v���7�����K�yz�MdHIa!�����>�,%����(�h�-	�0�qH-���އ����͗�j��6��ą�6cHYG�������o�S��Z��Ѓ�͝����q�}���\5%��0\�K��冢�3�Έz!���8n�`�M���m�I,�T�o�D�]ņ-��aQ���f_�	�.��dQ�1\����j�o�H����-��uХ�y٠o�0*)j���i�1di��7�z���� ��5�J�Ȕ��iU��o�JE~��%@GkB�/Y��1T���5��u�@�$��b{��yQ���]%1����&dRc�����6L�Rh�4���{y��X��vNI2��s�$�y2�j06�l�Y�"���R>(��{{V�$$�b�fD?/̦d��Ot툰./.4���Z�@��J��rkN�s�oI-)�KƷ֊/�u�$�97|� �ޛ\�@����g�!���P��a���97�(�e"�3Qrly�O5�׉�\�3�+�q~x���= �� e��j��p�OX1��:Q=>����=�5d�sIh}���K�,q�@�_zo�s2��?��7���p���KL�w����c�� :l���|� ��/��R�_��!�A��y)��^��z${?5@
��Yc�r���7^��#��1�0p�J��:st����:�s�-*I��KkJDO?;���D^�~S13,h�4$�-��o���%�;��R��������`��
S�#��*��<;Lۗ/��kWnfw�Juﶌ��L
*���n"C�}&8:���y==�3^B֏ٔg,N�M�j�ꟴ��y� ɢ�kR�xe㩅~�aҔ4�n��EŃ
����pr�s���I&��sZ�q�6q�[J�>Bp5o���D1=ҍ����~�$�Wa�\�R&{����-`#���p�_�a�6�KW'�Պhu���$.�?�MpaB��W"PkT=�|&}��.�sT�g�Ւk㖲���=#@�x�׆��p>�"��QG��·���	�I�G#7��i�@�./V�'��$�=j��Ԫ�����n���B����`�ph�%R�h-���X��#Hl#(;:&k���98��Z�_��:����C4/��	��ng��<���\�[`��������/�sC��iAy�@l����1����'�e׈��o�f��������6g�(8n�����0,2]_�"Z5v.���Qu���A#2���ѻ+pWvF6�O3�<]�O��	ׄ�*�<	@��a��}��&��{(92?�t}�x�	�e�0�q�gM(]	o�����-�5�SG�\p�T�h56ށ�>�<|�ФsGP��$��J��7� ���A���ʢ��p�����U7s?���M��LO������-��B�R
�jh�Yִ���7U���_/��=eF���g�9+�/���ERם���������1_r�;@gƓz�6����~���3'�R�gv��Jo���p@+4���b�54�{U?��[�T��]
�
�/&3��C��q��kry�%X���Nv��Pi8��t2x�xG�A�B��!�E��MࣱF^��\Xca#��ܯgF�ޓv4D�Q�L�6�a�Ο\k�N:�����95Zil�F�+�oP��Q����2�����ZI����D .d���ő�
/���g��5��Z�w�c�Y,��:�=ԯ�n����0#�ؤo[=܈�$�	�*��y�����ɧf����Qü��e���2J+�v�Ϧk�z��5�2 ��ON�7`>&)� �#?�ZdL�]�H���BO��҃%Z����VZ9�~y�-�vG��|��a��g�����
8kf�G������S��0�b���!�+���J/$H�@%�$^:�O�1���߼��d���G���������;�z������P�����(A���o�;ؒ �(�{`/_A�Np@�4Vb�z�[V2
��0�F�s̥� ���`r�#u�N�Vepؒ�3��W��Ym�'�©��>��Й(}�A�Z�a��|�u�a��b�h�c^�3�N �6��S �E#��BL@�g&[?iY���6m��Uӯ�d�W��2W7�X3|�����7�i��sM_z�E�x��Ȧ�1�����5L�HyN�e�Lh��:m���vW��Ր���;�t��!���Tԟ�L?c�+�I����#�5(�FCnQ|�Ԭ�w��Z��(f����(%䁎=��%�A;�ki��=�����x�Y�_�pO��u�>��aiʪͻ�v2
C�3S�%�����t�5*����4�Pz|s0��o����:��ի��Z���-�^��REM"&H��}�e���ć&�}l}�^.��D����1� ўr3[*�FV?Հ��	T -�o�xϹǫD�3y�O���4e�4mv_��8�'ݤ�n��/\��f��&�S�m`c�]�#]�m�@@�m!w���`��&c�7X��M��$Pv���L�¦����뾨M�]{�ɜ7��'�r%��/�{�6�K�9 �xl�e�J���'�sR;j��Y�g��M��6E�ШŻ<dJ�eOi���RO��Ӭ�J��L�D��%h�EH��˽QF4랒.�S3��<��8�g���ԼiiX`Vo���]Z�2U���;��n�;ؽ�>�.�xYI׌Zl�g=�h(���r�k|��1^�b���cT�����^����_+�,$��AHt94KH���z���3}����eh�S��Ɛ�Btr^xi����}�����񒌴
��/ﻀ���7��0�(Q��U�M�a?���5 �{ =_/��o�Ä�Pa�b�;��&/[�������!c��)�?Ku����./�	>�E�|p.H6(��Kj�!W�@!4d��nH_��h�j;>���Qxr"*dz&�/2K6L����U�d�>�'=f�Y�lY�<m���+��^3��8�m�f���^-Lǰ�Qb;�H�J��ӥ����/����@@����-N#B�`,o����FĤv����P@�0AH��)�
�)'Um{];��=�SRJm���\ǔ%��,�#͝��jaĭ�`2�����u��@��t8� �S�P �v�n�d��|�g��x��~0�733�G7�����u�d�{.I�����S�:�эI���:	g^�N��t�/�aO�lL�q�>&�07�
�(&�]��iL���m��b�����^uF��T��V���n�����&�ݏȁ�W���F~��e��`�]���z_vID��H`���1C�慫&�GŖ,[ �֧\Qt�Nm���Z����`(g�v�NvJ�Z�9����iXlxVHYEB    7288     570F�/A,�X1 "Cv��鋋O��x&LX����N��LY����QH�m=�c~I�3	�W*�G?]�a��e]w�*h��7��-"M?u!��@��x�Y;k0�Q����]o��=r����yҾ�i�JhZ����eXƶL��"��㏔jGܧ�O\���{�����u�n��h���r���@�|e��m�)�F�K�?�T
]�9�d�
w�ܘjʹ�u�솬 iV|��mk6���S}��7^��o�P���9>��u%�cE�(���k�G���L>9�z�׬R1'?X5�a(����,�@��~{� ����a���Nw9l@}S �؟��xU�eu)����y1�N����p� ?$%�cb�Bj��̉/��B�)���퓋ܰ[��9���}��0����?��:��4~>%��g%@�B�K���v�ܫER���F^�O���b���:k����B�2�	*�.iC\������A'�N#T���/${�-�FF�M&�c�}����,�
{X�C8������(��s�N���y@N!G�Fq�Kz�/T���'tlwA�I��!v$���z���2�t��&8�.K�ii܈�����K�X����X/��	�(�V��[��������(n�֮��#�=2� m�H�S�rs��V_�$�~ڙ������J5;my{T�FFV)���ܙ^Ŵ��DgzU����_󦋔�M_��5�ڥ����6��C�O�������櫃5/������ۖZ��틒�11�w�M-�*�e�YJ��i�y�,���S5�t�R�maW 39��+QX}�w��P��Wä��L�D�.����⤤=�iq�4��T>��~��4�t���X�koĔ����tf����+�>~	F�:�E��Ov�-0n���� �}��_��3����N��	��;�i^���@�cE^�jY̣�����i������b��ؕȷJ����lSDK�R۲�t�����E�*nF4-��hA8�K�]i�3��x�디a���
o�נXU;ڀE� ��M�r���*�mn$8�Ϊ�eD������K-��O
�Fw�M\W��;+k9�����(Q�іxb�ֶ���@`8�?��U0�( ����ܫ�,�H~(���,O&�f�����MqٌDqQ���xu���03�{���w��{��iԐ5Y��ۆ�/v!�AX�o��*w ���Z/��3��$b�nkRR�h
�Ou���� ��9.�}:I
b����O:�U�c�2ř���n� [OUŹ4c��h��?#O���k=8]�NC��Ve~؉���^��j�6��|�[=��9��b��bC��m