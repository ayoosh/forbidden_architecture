XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����l�T4$�h|\���v)��,8��U'��M�����nu0�#�[��1�54�>4P�h6@3���-֞��W�ع'j}�������v��_۳H`�P�� �y���z�@R�[Ā]}���dv����@'3�Lr�.�y`�� ��
�Hb�5��`����P��E�iѤ?���U��,�ɰbi�ց��f�bpH۰2a����|�g󤻎Ja�� v�P)Le�oԌG�j<ݐ�e�]7>�Fc����-N�..�	!�D�ƃ�~��d.V�1*��N��G!'����-����w���h���0C~���_��;I:U!�����y��t���cޚ�Q���YsX�4w�\�)U���_a������3z$Գӣ�������w��s,�,�b.��$���Z�����h�IgN^�s�"FZ\�����wWmMӭ������x��J��/���l9T�n�u6Xs	,y�W�R�)�͆�m��~���`ɐ�k�DZ������Z�5��s�=p3t�`d� w�e�p��;n)�%��o�n+�O�*��m�n�03ONp�q�3{@��I.��2�]
�pX�M&�]�^%���/�6��2�;�_+A�*d�S��4�FhH������l��~��������F��J��,섖�$���@�U���!}��_�s縍Ew���
�vc�m'�|^��X�ڳ�9R�����}�ϲA�*�����^��]�U��;���U���Xd�璪9��~_�����V�-XlxVHYEB    fa00    28d0�[�N��>���$o��6��mre��"���Wt���͖�0HB����O��'�HZ�4�\��'�C�Z�{OX�R�mֶO�j��'��=Ӏ��U�!%���~��MJ���qu�� ��^��Z�t)��-�����4�kX+a������1�gLX�fv97mw�x� h�꼱���:'��h����O!
M������(eTESR�!��*�n�X��{;[떃�wSC��� '�U;F1m�ӬcE�
K�:W�K�vD�3^]��X�|��S��w����+=��	�?�ޟjeI�5�MU9��݁o;1u�t=4�m�N��ծ���v��'J\��ͬN_�:O�G���䱎h����\)os��6zE,4��ݖ7.�����+��v5�2R��9�h�g����/B�O������8�1��wT[!�Fy�z�>#'��׏8)��9�R�+����`=��Υ�Ӱ���?oN�̮c�\�'y!`�"%e�"ҫ���R������5~�_���U�b�Sk��H�3l�"ߦұ�L��y���n�q�ϼl�*�%:н�o�@cxGd����Z��0�RE[� �h@/.���^���:�J�.�)�fΈbw������%1R���E`�Za�o�_����Nfy��D
���eMu&K�1,~)h۪���Ґ������5ڒ����8Ѻ@f�Dg$�g��F����WekQ.���*w�.�k��	�NZm�ڈ���k�r6�M�b��݋c'1�:��"�KR�⊏2<�޳�����|��;C'Fᔭ���¦��%���T��JA~�?'��ZJ?�P�1c���?�����%����* ��)l�\p��V��(kӉ��w���#�1��'ȿ�C~*G翦g!^�EV�\����8�L2���)���;S��Z�O����FQ$� ��r�c��(���y����Y�b߰kJ����mp[�F�s�<Z��O�x������s�í4),
��k����s(��r�+�nl�Ш�H��5�1kv=��pF/����^�_~��v!��=�$dq(�N�Ҥ~����F7Ǻp��f]�zWd�ؕ"����s��W�.�Oe	�T:U�CJ�[���8N?i�����F�ͥ����׬T���qj��[���0��Do�VX�U�0���c�I� ��N���CL�rIdǦ�)�Ϙ+m⭨�Xܛ��@<z�M(�vR`-j�������V��@a.��j��M����S�K��MT51�u�vg�,�@�ڋ��$���Ƶ��'�F��]����*B��o�p��NR~n;�m�}"	�]@T�R��7����J���GH_��lOe �H8�JQ���f.y��:��x8m�OC��ѵ�	ճ}���ܢ߳HfҔ�0`[�\��˔獁V�ܲ�ـ�{ԁ֓2�{�:Lh'��H�)'h�߈]����j�6-�̤�f�®"���Η��|̡����J
��k�-S;R^��:�-��-d�	�⼰��V���q�5&����i��4���֞.�0��[��{����6�
9��0��`�4Oٌ�Q�h���(�b�����h�~�Z�1����~ל��Q�Ђ|j���gB��FC^��)ƭ�S,�{N��e	y���MTs]a�.-αI=��A�7 �Z��B\s8���^��U���ɪ�y�RY*&`37��N�w����V̂�\hW���f���h%}�Mjȸ�S��n674���D|�-���l�����]��œ�w�G��_�2��v��vK���J���==��hu���m(�#��!&q:[�� p�'�5��qSh���Q�W�ee}]��=�\�r����s�Rv�w�S����r����4dl�$rR�T(���Ҧ��0��(&�4"�븊��Ae�`�ܢ�闆G�%Q܈�cN)Um�]�kj���uA�����qY�]����-qA�2���ʀ�-6�^�Wdʧ&�&&ȐI�1��3��������LJ��e�5W�4�
����(s�6>p�.708���2����V��S!�Q���C+y���k#f�\Ա!��5M$�����3c�)4�E	�\rpuXA�Å�ֻ/���aX�r/�hŊQ�a;{��c�f!�B�+�X椟��!������k;�}��^I�����y�u˯�Ms�o	t��*=��3>�˗�w¤����^²J�b>?�&5��d�ss��	���V�O,Ix��7ߞ&C�~����H��x_Ps��!����0+dz:P �j< $��^��?�7{�?ܨ��A�v����B��
G˔W��<��q�y���$}�-خ|/s����sBZ�/{�Ȱ��t�xX�������~9�Ü��,�K�����/'&�q���~�e͝��	�91�^��R!.�F:*+�����܉ZKAV-��*��,����Lq5�ɑ�U
����j���-�`^���Cf\u�u"�ymv���o��@,����M]���~7אɃ��T!��!������9�2�Ϫ�Os��|�-0�MU6ɉzq��à=An&���dޫp �5��HU�+�[�0|�fS X�R6�q�-.���e;���A`����/#Qk(�W��oy��y{r՛'xr;)�0rO��Ӹx��C��L�Eo;���9-�2t�b�ǐ����1�
?�&����"/=xk �4 �s��ɇ�o^j�:����F�;~��|��f'[�[ ��/'�!� ��yl4�tck ���>���G�g��#D*pґ��Rz�y�Q��!�
��`�ɭ��>��
�[��̔E�%�&�N��]i`7�xe%���S0�y��W{���m�Ά�ф�����90��Ny�'�����_��%r�)McW����}�f����)?�
��Y�#��(�)�#"�M�^dk	R{��4U���mZ1�7[��crׁ���{�{��K.9�ǫ��V��牑�QV2�ȧ�LJ��ݎ�n �V~s^S���������{�7�qŎkeBm,&�2I��4�ȨoZ�핤sN�(�$��UJA��KT��ݪQ�AK0)~}�{6���=V��"Z"B��䰕�f��)�^�	ۇ�W�b�f�
�ǅ�XmnHB.'c )��FBj5O�ڹ�n�M�,6�ǀ��j���/}2�_�����n��S�jJ��5=޼{xw��bKw�������i-�2_kH�i��ut�S�Z(jb�Z��h��g�����N(� G4���z샘{b��٨��P������E���c�H����nE'�����-P+�����&G#)d�*\���������k�+�S&!�v�l��S�'v
@�����X��HS)���t�j��s�Ӿѡ�5�]E�KjnZ���t�Gyw��a��%h/�=^��@�:�����g���h����rO畞耲��/Үk��fF�AT��-Y�2^�`�W�R��5�^(/��z��w�P�;Ӿ�������)�Q� ����Y��!�F��i�}����?"(�\ߑ�*6��4(��e�1�fO�+��L*��*�p���VۑS�2/�x0��*�(�� /'���A�> �y��P'�<�mS1�}�^4������>l+���∲��8u<�5����Ivnގ�K���r�vb�w����)6O�`��y/���v��*qc8�7<�>hM�m����Z�ΧV�)����T��9�9�I�`�Z��8 g��1�����g���/υ}�4]!1>�Tv��Σ��J��r�Jn���T��N
p�7�ː��a�X�3Dd����^LG�y���tSQg��
���q���D�+�
�m��`>@k|_1���t�]D-\��|:���B��Zp�4����ب�yr��N�Q�T�Q�����Уkx���9g�nl������ܒ�]�����/V��-��O��',�eX�}y�݁ò��Z�L��^ߗ������1||�ˁ��DS�7Ll��9V��X� ���5�(i�3��~�2���J&���ܡDVC#Y)�~�iϝ��9z�����V� TżQntu��'��bⷥ��ls��#5���wX~m��Z���悰�l�r����T��><�cՎeQٲ.����(U͗��e��I~$|_@]��G}-��*Tb@`�	�����5�6f��e��Ks|�vl�����H�*�)��j���X�p���(aS�����uLfA���ay<��F+��D�1�q0���� ���a�4�>R,�'x�����y3�Dw����<��	���|.�(�����bԇ�@��l�'(l�̏���!
�G#`�F��~D3�R��زW��նH}�+�p߂���Bo�+��x�}WW�"'i��T�EY�<	*Z����r���� �?�A�����7�==��aG'5�P�����!I.}`���"�P���Tۜ�~�ER#�4���ᓅ�O��89�x �"���x���g�%��ҥ�&�������`�'�f���,�?#��2a�Q�yG�q�u���Ѻ@E�DQ��x�KB�����
sF�����x���g�-�D0�9��J8�t����L>ZUM��+�E-N�;�N��db�����54=o�s��k4M�\	8�-�[8�^D��+�Z�7�D�@��7��)���>�
o@#@6�~P� �l��y��5����u{�,w���H<�z��v"[�B�i���&�o�\�y��|����Z>}�!q�Z�-�u�4�%N��8�������!-w�Y���n��p�2r�C���zb��T����6�:�\�ϣk�25���E׿��	q��kM�x0_����h>��N^����>�'�a9�`�yց��-q�5�u)O��$ǘI�Ė��#�G�8����t�=(�v�|���`zs����(�F��:#����H�l!�2:S�k� (	�/�L3��K^�Dh)�\�nɋ����_M�9�n��H6�/�[!q� �.�q�����n)Fo���%��9!���x+�\��$2s9oK��I�Ň���_���!��da��I���TQ���"������?��)9�$���q��+b[cQt�5	�QY�P�cOLVu�Mu�s�* �[���������
n��Y�{���uX�@g��X�]�Y��+H%�����>�O�ϛ;jQs x��%�,�5��;f�_^�۟ߵxa�N��pB�_��W+R��F�X�
�i�"�tt6��C�>ӎ]���V�*!KCo����W^|>v[�nj���6ɖ���;� �g�Z�����ݮ�����>eyPj�R��L�/�xђj�iV�wA��}@�"~4hFc�vD@�6.D����_{o��`�5���;��oe��U��'���ńet�U��+�����/�B�:��%θ��������A?օ��lBK�/��h0<�`�f���P�C��>r�����@"���g��%�R��B��;.��U�Q;6�RU�-����k��ށ'� iB8������;��ޣ����V���@v���sj��zqٲQ �9[�U�n�ݛ7�K�5��m���-���C���HX���r��I���V5�Z6�TSg%n���hU���Nq�|E�u��x�<��`-m"��ά�h��;Ӫ|ұK��
���BFeA,T�5S����lV���
"D��h����Z����};�͈�(�؉w�-ޛK������4ΝI
��g���)�����e����#��ț���oHt@���/'�e�0��
`s~Q�����ZGA�qO9�"V�0� ėyÄW=���\-�����4,�S�q���__ن?�E����X��hZ�z�8W���'�1]	�2AI��Gq�3,�5��)�7@���7�wrV/<�7�_-�B�y�8��C�mD*��vdy�Ȁc!��X�b�/UJ4=����aQHh�ʓ����ʥ�8��ǌ;�)z*�Wk�	��w�lO�j�]��U�U>�b�+̉U���n64���$d�% ��Naj������<��M,�9U��F���12*�L ���j�F/���v�e}�����T������
�ڼ��qU�;����)�Ni�qÐ@�X���(߀�"VѼ(�H���8w�Y�J����Й���W��`�2�}�����E�a��)bb�/��1pf�?㨂%�\j��w'ˍ{]�:����G���^.�Z����~��}�@*.�8�6b]T�6��Y��T���=s�Ӧ�ޅ�$�S� ,�%m�-t
�VV�tkǤ��2�Z@zl�I*�]�&���&_�=��樜�Q�y�0���+ʡ|Y��S�X����#]_,y���]%yn/�����_n�4T�����:ÿ�M�ۓH�tJLJ�-j�WH�x8�
Y���]�Y�&�=��,��/�l|c8�	��\#����3��^�-����Wl��q&u���`{�:�\�"q���֚\�cW�u�C"�t��s6�3�B�d��~L\V}q���xnGPp  ��u��LH�vP\@d��zWy��RU�X�?��+QP��$�q`p�%�����w�>�����-��;5=�\:k��Q ;I�P���(*��[y���sr�`�>�8|��hb��߿јSjN\E��5���0%�q�6D�p1���l��Dd8ϢvԘP�*�W��ŏ�e[VQ�D�X��Q��ۈ�6q埝׭����f��l}�4O�U|�d�����{_A/��ayP��+���.�C��椶�U��ghP�_�Q\7;b	�+�5���������$h�(��uq��o���?�螲l$⍷�=׸E���9�a%��w�dwTc���V�7<�I�֭`�+"s\�ϟ��܂ ��iGMW���4��ˬ��>]�\|y�!䲉v� 4�BCȯԵ�'����J&i�]�#�
��ͻ�$�Z�&Ґ\�R�Zx'@�����d�j��k0��VyK?�χ|��vՏ��pm��	�IX,���Bc4'��b�KuQW*u�j��l��ƺ�~m`8\���g����.j�@V��pB��B�;v<e(���4��ւ��{CT7ǲ�|𭦵%��[��l�� !יw�x��h~ɭ��L�𯆧@�����r$��B���ٿZ�&��pH�W� Gљ��`$a`��D�}擞��p\�e(��J�a�
��n^s�c%!H����Mo�,�\�a����J�2,����`qv<�,�%�Wc�6�Qמd�����h"1|��1ǀ�a����~	�ˣ�p�E7<���9~LJ�ڴ�����U��	�`��B{���]m%U�����O��ݽ"V�,Yv*PDs�jW)P�g��T<�F��*f"Z���<�_�����}���9��N쩟��齒�*�cM����+�	t��=�J�����d�f�^5�`���@�ȟ�j��\�u���\|����	��x�T�n��9��2���#�I��#ş/N^S�(q;��C�c��P�+�h��1C�:���q���nʓKR汔�Cp$�=�s_�6n�I�Dg�
-IO�'	���1Q\�~���X�>t���2�H��� O�O£$��Ц�:B�Ų����|�R�kT���8(w�_��)�\�FE�� '��T��^�M�CG��z����nan������_��b:t�+�ל���o�)�N��̍�@���U��-h�3�6��1�u�=T���m���	MV��h����C�����z��� ��j=H(�a�TsŜz��I�x�r�Kg������}��pع6tv*e��� y�зV9>�`k���P�<�>b ���?��(iɃǪO�T»J`��Jc�W��#
��=�;���v��H,%6M+���"%����;b7�����U*9D3Oq��^�я�cw��v�c���W�{Ӵ�h�t�<���{E&ב�Ѭ��1�R0���@���R\�����Յ7�f��`F�(e.)���t�/)N�G��_0fZ2*-�����1qi�h�¶r7������;-���Ľ�ej�F�2�����a�}��s�^��~�ɮE�	�3ԌR{�24~E����ӘЏ{��ga�y<����3���{��[��F+������xݛU[/A����3-�
?l�kj�W�,O\��~P�-�L%���q|gf���"�<}Jŏ���#I��G����[z�}�8p�{¸]��c�4��u�nG��k���l��'�|R-9��x߁����O+���I,DܴC
M��2y�M
�U�z�Ҍv����A]�g����|�V�4���X�cx��:�1�.��v�>�����;��I x�͊��%�v�Ę+��.@{���^0�(�&8&ѓv��;�NG��U�%��i�S��r:�-p�.�Ԝn�߶,ݝS�1�h�^?�S?|%���\��SV�<_`�r��H�8ԟJ�Q��j������}�rc�os2CWMƺ2̢���>����yr��/�۾눻��<���
�j2��ۆ���*]T
�o����'�^�-I6�>��c:ótuҬ�O�r�62F�����T`���T�zF�:Pz2�
����W��=��iXC��P2���/���1������H�4u��=�
,�c
�cA�ru&yR�����8E�̵��lY3�Pf�%q���UcΘ�
/�a�~�N�Q��l��t����<X���m\O���@9挨�Z��W�N��R�U��}g�,��^�$c�@��A���o"�y���Իrm9��\�m��j!Rr��<��%��{���DCZ����o�`^�lGvd����g��C'����C��µ�	��i�4�ȰzN�,L���Į9�aŜ�Bp�`�����}4���V�cp.E�v��}E���w�s��74;��ˀ��v���XN�fX�@���.������be.�9	�P"g9�ju�,nw͂� +Sgr4<���7�OQdݓ[3�ϼ�9�I�GG�x@��AS����.N\��<3+�S��X��{4@���tj�d��Ȩ�S��"}���S���73R��o=����ǈ����t�# �F���гG�����P�uqC<�b�LL�����a���:C����}-[_^��@��":�Ɩ�G�@(�0ֿ�v��|�*����!�Ɣ�����Gҏ����L�i(�߈��z�Z���HABGix����?�
��"�p?�{��7�?����ּ3��$)�(�|�c���?����9I�� �h���:�QE�X(7�IRoT�N�U� ��(�l��w����,��9%���u��H�N��&Q]~��^J�}��5)g.��h���ovOvN���
ޒ*;h��^��"�4rELZs���4�2�&��(B	���oCm�<ve���4�k���8�yU�Utҿ�L�;x�_�5����9�V1���N�+��q�nƽ/���7�f�H3��{�p(���"]PnU�)}]k��^J��f���}V�n�U^Y��r/|w�b�db�+��� �+�S���s�8���b�M7b������F3�ɨSj �H5�ce��'	~$k�1�w���ĝ����[��������f�[�/I��".*����p���9ö�;ґ�*6p^T�:�W�B��/(A'9�����&{b��鉖�������jy�jH��X{�(��4����b��Mw3�[�z� K�Dn�?���&u�6�	`��L��g�w�HH��<�������̈w��8���%D�O-���۟�i����꾩�ـz�C��.� ��V�z�%ܩ2��E]�R���:��%xm/�r�ǀi3�֝A�E}G�`ҿ�\�꾑٤Y�m��o].�tF�Aw�mg�s��c9�7�/��t��n�V�ʄ����@�fwXI��lV$#� +�t2_�9g�m���C!���6��@���Z_3zR�^���0��HN�y��<{r��^��T�cT3��i����S��9H������#>�=>Zu?����'VP�w�ַ=�Zl�aX��#~�V������� �p�CܿEQ���������gS��"ֶr[����,dr\�z��b��k;�C�
h��L'1�ҠL����>�O����]|��� ���OXlxVHYEB    5f88     f30���N��B���)�Pƻb�0!
�q͋S�nJ��-��+�A(�x9�Y�@�CU�I��A�5���5�D�(
�2�,��i�S�p��e�H�1��2�ǣ� ���QD�/��븐�,x΅Q��Ѧ�5�M3����[�,}�#�[2�"A�5��ʜP�ֽj����,�љ*#.AOj�uO0���^�g���u�a��$��ZY�
�ҋ��q��C<*���B>36�.^<9�	P�'��b���L��ɢB־�bƹ]4�fɼkhN��Y�3�P�R�W�=;���%����fy��cd��NQ���|���w��p���#��;��7��v���_`�'/w3�S�'��n|��Tlą��� �T����'8c�>T4�<�%{����Jz��`��Y3�lG��޵����[��~݊^�?�3#���+�o�g��ii�c��e�sd�ZB�^��`����T1��7V/RU�t���s�
~�:9����.��9�@A��x�BOB3��)؃�V�N�T��"��������1��e��]��8�:�S~��@7{�V�ե�� �do%=��M&������	��ł|��(�/������]�?Ƈ�7�t��Ev-��Wq��?o�>��f����f)����E��N�`�)Ʉ���)�wh��vI	
jC��Q��A)�o'�j�?��"hq����@��(U�&ho���s-��TĨ��������H��wJ�a��q:�MK`�ꪢ'K`�������O-�$_*A�%^r��D��-CG��<S<�w�M�m���]N���$�x)���̢Ef�)�����6% яօn�1.Xa�I�0�7�I�C��y���S�omךi�:@,2��5]莎t���t8	�(3;���1��a�$��ZI���[f��nG��N�� ���K,$C�$�Z�DW�)z�z�����}{ؘ[� ޯ넽^������?ol�U�����<�h̦qP�U���3��`^؊ּ>�cH84�a�����{�ׂҒ(^����}��rb�(��(�9~M�Ii�޳e{y}��(�+�8|+Y,�	H0��j8�T������+Z=|��y��'Cb��҅��,�y�b	����@��b*��-��W����qv?�?���V��XG������h��rƍ�c��Cf�Z�Tq}�{I;�/���$YhK"�"t��-������!��N�lg|{5`޹;����9щn���<�j���u�;8��	��7�ѩD��$Qe��˘/�~u	�Y����a�?�����%6��[q����{�����+����1���#��o�<�K����!�PW�vW�d�P��Tcwo%�䮺����K��J>g��W.�5@�7?�1�{��/��~8����WKI{�����_;����W�I�,�\��i,��"B�
�[���і��4���F�wbqވ��7��̻yh�9��b)�+5�r4u9	��ӕ����|쎍��g����6�����;y�5�zW��RT���g@e&r{z1��ڱ��L�A���&!���h��������,q.ۛ]pʄU���!�^�I����.#̌�M� (<)#\�%�c��{�d�^O�Jz�P'
2t;���T�=��T�=��x�Uj%Ro2ƹ�:my�	���`.J=�>C���t�Ө�;#G*��_Pz%�pM��J�-�R�A�Ɏ4fXduֈ��}�-��2�\��
��I���&]�x?$�.�	��܃R�2�x9,��8BV�&���j�8��Ga��t:y�(�������5yG��v��@�l־�0J�#���?�v�[ő)�C�hA8���(�|n�Y51V�w�×��qn����;Gb�*1���0�l4aD��'�A:��D�Hjd�e�ޮ�%���ʍ�$l8ϙ����yq�;��1�E~9h���BD�広��s���͸?ػ��mG�����5l�b�ש�ކ�x���h��_N|��SЭėՁ�T��/�������0�жa{�P��4wi�%ȼV9����Y'(�i��0�oP���7��>�<�SL'2y ����z�;��?P��5"_����1�YHSC�S!�v	��� ��r!��4ݞ��m�u�[��6Ҕݔ��2y� ���r5�]�1��R���_\���-�[�;44�*q�@��Q��1>��Kn���Z�Σ��W�|)d`p�{3�0ҽ"����U.�j.��A�^Z:@Uဃ���m`��+�}KCӺc�G'״'�:�B�o|����]4u~єB@��O�d�͏�x]N�v�5p����-�[�Z*P��K^��X��T<��	�O�%��ow!��_���;(����
�
V��R5 ϊ��k���iC�E#k�-I�3ۉ���ȳ���|����q/�y-R������ c$_$�!7 ���J�����!j��Fe-(����
����/������%�+v���I��ԋ,4\V~�4���x�C��r�^��M��^�6�m:�4o��K�{�N�/���P�W%�p) �ZN�!�.}�J�:X'<��i[�*��?���]턑̉���@�d^=|�~��][��O���+��"���~;�ҤΆ�Y��me��&�jqT��8.��> g���X���j�ԓ�|���K�!s��kٓT��k�W.aMM��P��o���4����V�	s��Qa�.�^p�!ha�,uu���v�E����=�g�/.d2ˣ�N��uhrdyڀ&�<`�
gϦ4�gg�5NUh.��z���p��qFP쒴S�:��E6"��&���&��
U��<��㮕�ps>��X���y���5O�ZH��[���
1����->�u��(���M���k�E�4�G�uD�[
n����&�g��]�02��_�F�1���B�q��F�Oz��C�cB.��#囯.�V�Sw����yg��`4m0J=�]ť�'ka�N��i�U�K�%�B����UN�q$�\�F(7Xj�	��,��\Т�͕�{'֖5��kX���� �}�p0*�''�%]CI^��0W�uLê�{�t��/�§+���2�9�����¹͖���d��"�"�+�?�d��g�C���N`�	�pw��~47>5=rh�3U,��oF�,�2�9�������J�n����l���!AN�ծ��G��n	�)�ɲ񒔂ɴ,�o��O�	��]�T�K�U�0p�t�F�F��t3�Rs,gP�Y�a-23��7���q���ͽ��)L���Hu����$����;F��ۅ3/R�_~�!�`?���L\D]a_�z���&p�*-�K���.�]5�E��'��q��RBug⋎I�ۓ���,��xW��ڤ���.y�O 9��Q1� �z#�]�<�@(\�.A1w@v�Q�n�� ����|�f������� l�m�+ł�(��gf�=��3v�L�>�E��h�MF����Pg���@AG+g�Z�uST(;�pn��C��0����Zf���=���,���·y%^�('JP"i'�J�p���̀WԂ�C�w�@���X3)�EƟ�I��Ѹ;w�)��gT�֖
���|j��Z�[�=��U�s�J����ח�~e�10����Al ��g172s\���~�Ouq�'~�(��zy&���#N�uÛY:
����ϯ\67j
�/���@X��Fe��AI�Z$"8oYF��?�;m�R�������n�å��J����J�q��j��&���L��mݚ�ƦI޵:�]� _w4?�"v�ԛ��V���l�&lV1��J,�