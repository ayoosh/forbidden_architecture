XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ւd�� 9��ۗ�ajQ�!i��&5�s+�K�p�����W����!��f�u7Co���V��K� �9�P,y$���S��֮�#Jxd͞��S���pă@Va�̫6��O@*�H��.ADER�j�+��o�C���z�l�E���
7���LE�v��Fߢ�D�ŕ�A[1Z�������v�A�3g������H�,V+�79rb�AfFYe�H~5����i����$6&�˕�Φ�8�hʊ�ܺ�O34=fdV���Gk��r6�wc��ŕVN.�9���i�����씳�j:8<��f%3C�GW&�P�%�ta'�r��l�1b0'9q����*���a�;WH���m�t�<�XgC��{�#j�;�O�ڀ�g��?`���wAUL?�}���,^_W+|;婈����t3���sհ���G��~�E(��T�d�m��B4=dg�Ϯ[{����.�l�$L�B
�=wL���@|�'�k*�Ŝ=�xr|Q�6�U0�5��c#���T~�����K�3���Ec�����]�0�lm�*�U<��}/S��w�ś�q�'�׸$4c^���7��>���
�_	ڗ(�9�o3�����[��%�nf��C˻�9㹈߼�j����r�� ͉��:��d3gc�a7}K}wS�L:��b�&�]f�Y�o�A�ԍȳ�%J�q���)�X��$/�{���ل��(��y����7��~
.<�v$�H~����{@��XlxVHYEB    c67e    25d0 ��4/j���cI�O��Wr��}���J��|mN��	8�ƪ��t�9-9�v�C�y|s�*,�򤐧k�l��o��ĺT����hݢé�(����TS\X��Y�]ms�_��+�ANp�Ť�d���(�c�4C���ūX���3��N��k����[�<W;U|u��9�����M�2{�{�xX�%�S���䁵��!���lF��}7D�?�9�����JＤ�A	D(�;��3��� �����ɀ�ë���b���,#�^j���~ߚ�h�ai�����E��4��y���`އ��ӝ��݁ng��1^�R�}FT
�8�V���g�&5�*[K�V==M�����aC*%a����h��pj@凣,ɘ`�]��.��J��D�)o&6�dt1Q��CU��̷>>�;��~d;,�sY��6�[�z/)�N��o���{L�D��v�s]��8����U�β	g��\�A�*J�O���H���V�E�-L�L��."��e��>D�i�1�,L������9s�����y0���f�]Y̆�
�ƵSaAK�?�1܁x��yG�/u� ����"�$o�~�v��j����l�����ü��>��=�ӵ�6ñ�����6V���
fS$�ߴ ���
����^[�Ǒ���n��y��ˢ�@�$�B[�����ޫ'���R�l�T8����tjS*���t�A��.]��M_�y��~TE��F���<4?oF�3�"���w���n���ma?*ס5_��@D�#��s�w�_�gJ��|���\ǅ�b��Lvm�݃]�n��K&����,"�i\�d��@s�B+�WD\)]�煉�)`��Z�����n�6)��+�qQ�*"����벺��%�� ���+�k�|����<�u��vJ: ?��e%㼲�w^�&�x^)s_:+�nh 8�����	�p{�!�9~��>�0�v���p�ݵ?g%!��$We:�������3eD�T�����fqHɜnR�w4Ѽ�m���68 EvQ,�G�O�'��I>��Ħ�q���Մ��:'��O���e�a`9�Q�z�lNR���	���+�K�P�����V3�I��h7|v(v�9�K�!"P/Yge	��N"���i�QJ4�+=D����i�8�OWЄc6�	�i�X'����'���d$��	�xWa�E/
C��D�O���2p
�=��jT��Ҳ>��Cd8��N\�|��O�;Cd�PL���J�N�Ų����i]�����rA���A��|�,��,��(&	�:/��i�}���?�)�QJ,w cx�\�
"�u��&�����6Kb����+�j���g��@(m"�$�w�[h�&���o��]L8~<��K�z޻���z����+b��\wy{3%1ݻ��'�3�����o��Q�0em��?��'֚�Ѹ�
VH.0LV��]�V?ּ�^`�V_F������3 �X��y.l"�ދk �H	���v�����	��\B]�>�Y!VYj��H�z'���� ��c���hC�A��!`������0f���{N�����i��	����F��?���%9؀��e��[6]5��� ��B��@|-����9����,�E�U�z�n�s#�-��m|�T�C5�g|<qe i1�>�T�Z'�5�����thP*	�����-I��'L�U�F��A����ob1�dD���#YxͶ,�A'�򫭛qӘ�R�J�{�W��1�&�#�靗;dT���T�mo��k	�t�OI�M9��~�U�t~u�,�DP4zL�^j��}�$��f�²Y	Vz{◣�V���Q��I��g�KP�S`�ؓ�h��c |��*D8��v�B4�L�)�5}\�X�����}�ס�]���z)#���
S�]���p�sK�"p#���/����q!Dw�r�P�@���%�D�v�.z�"=����Z� ݒ�Ǖ�x��c�[x���[PNmX�[����)�	���Sc��z���g�$�P��a��*2ڱ�l����E�j6%�':10f�yx�+E� ���.<B��%+y�W����˳o}�]^��b>k ���1����\Mr)�IʍcNɑ����0��e� Z�Z����O���~�� �����㷣�$������4w*�@q���b�r6��u
��l�H�#��k�5y�`�8Do�]�wGBTE M>��#A����$y!��>1,O�7*1��Qi_{-���G��*|�L��U�4ř��qq[7��W�p�<����#�,�1*_�����V�V����Tn�s�
4��nڎ�)DUJ���%��#��,�FpV6�,�z{CM��M��Ph�o��T��/��R"7��5�P�%L�k�p*ڿ���k��u���]��&�0��_A��y�)�= qor��qp�^��#����*T�P�M��4�N7>��?Q�Z�q\z�B_�T���^�}P��_��u��R+R��)�v�\Vh��VZw�'Yq��"��cM�`�9���W��r����p���f�&Iu&Oe����F�Q� L���=�w�aKzۑa�4����wT�!��R����O��&A�B�Ψ�_=Y�w5�c ��~��9ހ�ȕ5�eET�:��w5[�k8/CX#ɚ��R�=$�z>������F� �����i!"ew�w��UN�f���3�.�9m�(��r���G]�[�!�|8 4���n�+w��c;NIG��� �f�ʑ�	�1T�;C���%�}WZ�p�0ښl�3'2���iqR�{�^�4��__��SP]NF�u
n�E��Ls׊,F	�#ҫz��`q�숉���6-�)4����ˈr�a��qlU�m'9n� ~:�2�ݥ�g@_�*��3S��?b���{���88fVa�Ks)F�4�Żf�5�
  �M������Ew����Z�:�Q1�q��f@ec�?��j �Nz#� O`�% >�����J9k�1%kZ��q���RYF�;��J~t�~��Q���H~7�Մ2���]�R�)K���X���Y����g<�чa�T�;T�O�Q�m�K��$h��J.=f�~B��@q��g��}��җ�##���`��J	�澻������r���T�ӛI�G2��{+�񊖣Y���[LJ��Zy����M������Z������rP��!Y�lo1�'q�#o��1��=��u~�3�_��tr��������M�!=�n�I�mlRQ�B�	��DRjso��|y�#Y?��{(l���i4��?6�.hW���	���Ԯ�U�Au�Y�Z�-�hܫ�b�(O��)$���4,YÃ�'��i�\>Bk6ؼpO����&�Y���|�~A��z��ǑDD�K)os����@��U��u�¢Ê���ɱi�j)(��1"����[�1�\��膉��ܟ2��� ��������x���rY+�����1o^��jڇ��>~���	���>�LP����^+�����q�xI�Ō����0rki�¿���@8.{i�]�����2�DD�����k��"��VBO�,�s��9=�7Z*(�ٝO5��P�������-��~�����Ҹ#�!�)����g.Mc3���=7Z�^�	�S
��"�5�e�Vt�=ADc��GEMϨ���_}�h���s7�8d§�y�tWo(��iM��)%������{���ӑ�5��."~_�<}��'1�L4�{*fZ��K$�jC�^�^ �[�S��ף7ʨ���H��M�2-#ኁ��T�ޞ�J7�u��a���^E�4v�^�2�	��@F��l���H9���ޭiTLH�W�\��ɱ$y�v7-h�q��m��ŜL���ٻz�����?�{�k"9jP�3�䐊A	�@�)����5[�D�CM3� 3�ԅ�i��}%�AEO{r�+��ʶ���c�#F�-E�f���c�X��K{�_x�^��/%Fm3�t����r�|�(�['I������$>�r�X��7��^��T�V��S�\���~M�ۈ��r�˩�W���+���c�\�paFc2�=v����h_�f�EǨRlJ�9�,��-*�E�X0R��/~�S���߷��� !Q�ʭ�+M��RKw�>G��-�4���b-܏N8.i�T��w��{ٷǑ�`�݋"��1;�mN0f�!��Fg@���mM�A �O��M<�k ]��h�e@��S���+���r�3���Pc��#B$c\Z7d�S��Y�У	�际SeH7�j��kd�ns���DA5�UE�
�T9M�P	�F�V~�V0�8ͩ5�;�X���h��d��h�ȇ�Mr�8#�0���_����ٔY��l���� �<;e�-#��e5CV�̌�#`�S��dTfx�&^HW�nJ%4b\n!I怖�:�*AM|��5 "�� 汕��x��U#)�~UV�#�b�L�C�0�h���B4sM�W���Jr�TE�f���֥6���:��X�\�f���³�>�=i�R ����@�M�H���d����h�HҼ��b�O�!h��Gn�4eC��K�Z���/�j7� J���ts,�\Kv�B�ۮ���sH����*���T��2ъ����et"5�f��kL��tx�\�;��E�
~R�Q���5��2�~���8��K�i6��j�g�	�e����]8�}G��)����e.��n��Mc�Z_���c�\�����9fl�<��*n/���*b����� t��O|�K�];����>�W$3[*�-�Yb��z�}_��N��I��^�8�_���_�0~EVߧ�Zib�Y8Ҟ[��<����݄��A�NA	�W��?%+�T6�m����sw)�{WZ�j���pB��ߴ��h�/3-��&}%`clLD��.�6r���`�� ��uD���ҵ��U[�[c�0���ț�&��I� ���K�G�o�'�-�i�Q��A�pҹ�F��3��L�L�`.{0Aѳ�%����f��-��YM΅UgY�A|ցXՅ3�熃ϣ}���N�I^��(ߝ�7��qs/=*�K�
��Jm�;�xKI&k���0oK���'6�dp��1��ϸ^ҵv���=$���Ԫk�ORj̈́��m�&w��r�֍@r�Lt��1
��8�t&����};Y�`Ċk��@����J<�E��lp���R�Y0�ٖ�-��0_�~�)]=��Ui:
+]�P��R��*�S\�I�WH����n�I"�^��Q�n7���h�p�t�\�-�9�7�Ny��?���b~oD�{``1Q����8a\��O�\��+�Yl����KT1�97�k��0�k����3ԣ���u4���7��q�^R/��3�Xq���Ƭ��]����*�St	?a��6�&����3C�6�e��H�� K�ϰl��3ݳK �O�N�p��ؤ�{�dEULr�0�,�A��A*쒏P*��H�V���t��5�Q���Wê�dl��Ɂ�(T=�� T�F�����@�!�7����*�-	�0�����`���2|�2�bx�5�b��=��X"u%����=��ё��^YOޞ=22(�蚤�7�;�[����.P�yyt��~dT���2pB\C
W_I�8A�H���n�լs�O���F#R?�l�:2�QiV���p�"Ͷ��΅��͈�q�W� �~|k׫�{�E�W��i��e��% �"9���D"ߜ8�tuP�g]�����`���7�ں�����UhB"O��S�����r�����su�>;���	���k��9BA��]�GrJ]{�!��FNJ�/;�Z���ung�s�d��0��:S*��5�I����$D�E�E ��I+���]ڵӌ�prvb�#)��N�����{Uk�בd�|�`�2:>�z2�<�]�'M��Xv́;njmjY;Iί��.T���������}�d�LR��	�1��H�U��TN�I<�L��+s��KY%E�-�{A�#����cӏlH�-鲝05�Ss���?��i�<�\��lY)J)��� T�ѣ�3�M�xa~ځ��������V� �� |
ӷ��p���9��9�r�?�W �`,��J	M���-���6��Ȉ2R�v��7IrLW�S#��e���	O���7z���=���\7�Gs���<W�lB�..��8���+��&��=�'�n����f��Kz�<hqD ��!��I\}��n|��h8�=�V�1O��g�ht>,ت7��M�PF�ׯ���O��?C|�RJYYj�Ѕù\ˉ���F�e B1Rl��L�3ú t�_D%�-Ē��l)��V�Ʒ0۫�N�II^q;���G:�O�������fp^��2d�|�a���7�\ӡ�Dܪl$����#�~6w����ˍ��)j�Cq����U,(���C)K�(3�E�'W{+�{ g�n�l��#gm�q�މb0��[>[c�����tXVO�z=�ĕi�hm�&���a�F��퐕����c_L��E��#e�,U٫�䫚��p�G�p!���\�:���
�c���8$Z�1u����0��וҖI�ް ��/Q�%�ņs�\��@0�������� U������#DeI����Z�g���n9���DN��kmA��1(SM~��a" ��'�����C���k2B��|�S;�������]��*2�#^�0�y��x�륺� %���d�L�#q��T�z�KUc����7�n�]N�Ox��;);���:��4��*�N
^4����-�g�ker��NPC�"|��ٛB�$0%څ"�@�M���q_�O�qӉ��U�e�~x�5�h���nc&J���Yr�o�W����@�9�u�&}���1%g�r3��|���yN`\ۢ˽�uPa�k=�^��-�T$�x@2�5��Ӫ.q�F�����5�׳���BA��֙�z?OC�#	�
:yz��H�`B��Nl<�@-u{�$j�v��,�z�xC'\�U���iC�u�o6�0l��ޡMy��0�C�rQ}��p��J1ůP|���5����\��5bd���� ��P���Z��8�-�m�3�@�DI��[䒤������� ��e�-IN֝��+U�I�J� �.`��#���QЏ�p����2���""u�$/xU���̋��ʞ����>\��&H�]�EQ����E�ʹ�V�$�N[���;Rm��DD0f鈿���S��)Ȼ�~��!w�u`XX����si.m��Y�p!X݂�Vae�<����"��U]\h�����ܑr-C����e�~Mpbje�:�`�	�±ڲً%4l���OH��M����o�鿛s�1A�;���G��`/%,-z� *6(��/���#w���]U=�oG����ς8j6T��M�2}]KW}d��:��Va����+ �\��Y�ɝ�� {Ŭ�@ٕ\A�}	�֚���9�W��ɶ��wܡ��)�Y�����(gI��X���3͌E<)��t8�6f��^<�D\r^���"�-R�f���I�+_rP�٘K3`ͻE�l�-��:tŖGynt��Ʋt��Ln�<��J�Xl^�^j�S�VF�rt"���Sc��y��;�����`ڈ�e��*��Uf�~�;�l��O�f76��d�ȁ���ʱ��;���3�,'��:T+=����U��j�UA_Y��V1Y�dDH�cja��ӓ�-��W_�r��㵤�ESh�A\�u����¥��Y��|���MoRdJ���	V�64�v������n�q�ֳ�����$Xѯe	=gP{��J�r��P���"3�S��F�E�]�9=�D����j��|B�L���3qڽHa���ţ���Qc4ӛ��*�[�^��<|U�5Ws2a1��4bd��w��3�����Gh�ܞ�s���Lv�v^�~��ad�5[��o���г���{���_�{��_��Ή��''+��@�p٨�92J5� �EFkTWL�ob�	9s�����γz�yw�(Ou��X��HA/��ڍ�7������Bv�����KLl�?;���B���ݏ���K���E$�*$6�"��z7N|��\֝�S��Ē1���ډ��Lu��U΃������]*WʠW�7%�ܴ����-�+_=�N����̃�2#53ކrɘ-I�J�Eq��nk���Emї+���ƍ6��9�� m�t��blh;���M��/�gf1���!���kptu�q���`���lSll&���)1+��~�-�f�n�}�e�-����4��>k����x�OB�A�Qjz+O�"���1��#)G*
�~i�%{�O�����(�Ü�I��K����Ŵ���'�Wq��@���9j�+����w6�����Y`G.���&����Y2��{��y��'��ɳj�.��|S��ō��(b�m�Z��h�Q��>jb�����8.�J��D�F�-#���LI}�c���#]͠�s/���@��}0HJ��8�I��9ǞY�􉜐��|.R8ri�)���/����r?�<�p�x���_ׯ��Ѹ����.`G�_���]�_v�+	��X��fY�
�pR��4*Pr��,��Cŧ�+���?��ű�����c6�%����h�9��D-(�߸	<�?�*퐀�ʘܜR&���;�@�+r�t��j,���Y����x~��M� T�`�4�C!�>�)��������ڵꊤBlcِσflz�^\�ڝ�5T%�������ʑxrz���P�=��T��T�[���+$R�@����W�o�B2[��9SN��'>Um��25{:���H�E�(`�H�{A,�Ktf�3����T�����p%j��|M�?�l��ΐ+���y�Y�B�j�ßvSUl���`�����J�Jl2w8⨇86�M�k^ͱ�%m�CBT�<�$�A��%�bj|�Ȁ���^�d�� ! |`k.)0�ة��x��]&!=>�Z=g��Z7�*�Y<-��Z�^�#���n˾e�O�U��+�ԧ�,�V�<��q�=��Nx��
�C|�,� *[��5�#;ӓ�f�s"�i/Ԕ��� ��tq���o��0h~�E5@8l0�D���C6_e����gb��*�(�X@�h��ٷ����}$%bE��݊��X��9J�gI���BR��mJ��	+(�3E�?f�)��@��W������^����u����ǧ�ه>�F58��iQA}˽|gQ�]4�������J� y9��
��9e��c0
鿦��{���@�:��� 1�Q�"p���i���
�wx0��럞�r5Fҷ�` �w�]��T>�"�<�-��i=~�[�N���%\b	�?@��[4hs�sF�žQ�!PԻϔ@y��H.�X�.��(���Զ���̙J8$ݔ�<�g^��_���G4��Wү2������ Aq��G����$HHB������
u��-�+�