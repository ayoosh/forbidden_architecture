XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����-�`F\e?�%&�/�|���B"; ��s#�KZ�])܇p�j�৭��;�;���=�D&������585�R1�$|��U%;/��kd�zB���%Fz#&�|"�+���afP�|�+�Y��)�D=
�\0��r��O�0���]��R���o�������D �WcA�r�gw�NJ�2b1�O�D��_���̓�kH~(�w�P���,vI�}2�-���B����_B��*?a��������Z�Q�}��.k��S^����Zѡ���+��T�(F�����߿J�A}�H@�Py�p�[g���*��gi|9>ȔI�2���0�Ǿ�-������y#:��0�"�|����������F��[z�W!#+�À4��� GY�{�JK�8�C�8�)�E����
�h�jj����.0�V���������@��NL�+�5���:}�7� �(��(~�|��Ӑ��{�����#�gA� �^_Dn���]�Ve[�Ĕ|�kS�C0嘷���b���}���2��8��_�7���ѥ�����=��@I.�]�e�PR�W�Avy�@�m�i]���#.b<�	����f#��朳�%��?;�P�>\���z4�����Cj�Yٴ]��'M� � ����Oi$�r������j~�+�ޯO�2B4y��.C:m�k���3Y��(^��'�r֫T��]|M��A2_؁��B���N����=�$	�% Uɇ)���I���6I�|KXlxVHYEB    2ddb     af0je�X.�7*'��!iw쨻�S�*$���HА��cH������]Y��71��|I#���wú�����F��9��A��B0�h��z`O-���d�Y��2����������2�h�od����Z�Dm��T^��g^R�Д X�a�)p'Ϧk��)��_�)������=���Rb4�>�~c9>7��y�M꿔V�B�2��%,��u��S���b�3�[�N��fXĠ��xh��>	d�,���Q=,��ā�ْ�`)OP��Z��[�uKY�QB��G�,��B�&!�9F7�9�#ο1��W�u��w�<�E�\��-D��
�~�A3�E�������IwEɋz�Ib.��QL�����]�P�?E
фo��?�������j�i�Fb���q�s�G�L�ܨ��/�y�΂_V�~O{�U��1c���l�84�~�P��z��Ch�3P$6�����C���g�Pb�Ԃΐ��yJ�0Ku����IE��x���
��v ���j����pR���;�1[��L+O+�����,a@�Y�u`|Ky�}D�h���lC!�6onʯ�y�A33u��*�`c�^:��CM��!�K1�w^�d�����9F�Jo��00�"�c����pʢHg��u���[I
����]uc!	�fG��r2�qD��R��6�_��j�`�?��'��я���jHL|�/�ݏ�ݯ�b�M��`&`�~��8~i���>:~/I� ����}T�[���y�fJ*�ٚY|7�!(��=��뉎%`�:�"
��.�s�m��`[<��,h� �����������V�/W(h&�՛�ڐ���RM�xtN��n�-���MX�uy�L���X��V�N:OI�ogd�mۈ�)gO~}C�-� �.c�X��I�pk�7�R&�j��g�,%`�>_*�E�"�6�U�}11�l�ĉη`�yc��RKn]���|I��6KS��Zr�y�����kg;��K�U����ݻj̸�d����I�ߑ�E��|�L����x�H �m�D	���n�w��<���Aq�3��9�.Ԥ���Ƶ&>��)��ZH�`��ލ��-(ꕚ��-wܼ��ٖ��o�(\Ϥg�I��J�0�	����Ȅ5��x��UR��yB���ɜc�E�>�hA$s׻7���=.p�AA�A�愳"�r�ҷr9+����h�:[`�2%��m���S�ax��K�DG��hR���zZ?=tU��6�3��ߔ�ʒ
���p�aTэ�Y�� [�|�w�DUx��ֵ�G$e�����W0X��GL�躻�}S�f������s��\���W&�C͚��l����v&|~U�lQm�wc�2��*���������?�g����=��b�U���$�2��X�c3Y�Ȉ*�{��+t����p�(hpA���i� L��6c,%ޔ��Z�����m����c0	㲖�	r��v�Q@�ܟ7:����	p�������U1��%g'ۓ��
>�М��\z��e߯�_��bǡ�OL�%�7�xh��^!����`�;�_�w7V$�S	�9-/�2&,�|�G���@|㵪�=��v�!A��	o �/j��-~$�Ȃ�Z�����7��Z|�Ō�|L�F�D̓�ӞlC�j�e��(�4���z�fk8��)sY
�1r����kv�����5/+�.�/���C�b(��af��o(��<c%��(�9j(�vd�,�ڷ�m�}� ��hz:�N֪"��ۜqa-ᦛ��OIϙS�J�g�P%v��j��������LѠʬ������tf�i�:⸥�����]�r6���E�?��T����D���E?8=ew�l�8����Ӂ_F%�0�%��~�����i�OO���1����r�M2��좠�bO�P'�%L����ּt��z:��@�dJɶ3��IkǙ�Ϗ	��F�N�^��5��0B`Pq~���q�
����r�~�y���L�`�Q�b���>>�P#��:�x�;G#_	{3J����?~��T�	ϝ�����Hi ΂Z�.��+}���z��0���BE�.���|M~JU�� ;��'r�c�Cc�F/��d}(��o�(H���xt��n6E��>���{��Q���*6�j���;����żzￂ�6ɊJ�S�НÊ��s>}0b�tdc��G{�ϣ�j���(`��><��IzS��)[N0(Vl�Z��U������"(�țP%<Lfǎ��丮]��e�*G0A�x��1��nWyls`K�GwA�w�n0�!��!��A�b��W����-��h�_!�����7�����S�2� ���
<J�DG�U�c�6�����ųn� ���W���Z'9�P��S4�b��;R%	�sF����W�3v28���wc^F�!S��䇬��o]8��]�Wo'�0��L�t�07�Q�}�"!�t�Iz50
�AU?����n��Z��Q,+D	TJj��Q��P1]:"�IÖ!�.M�f��zx_}�LO�u��/�e*�L���<Hɷuj��ƫ��՗dG���G��98V�E����Ȕ�������zY��Fmm;_⍁��k���M����}�|��8�ż�b����WTu��� ��m�L�r�)H�x잲h,|�aq=��D�-�,��X�.tu��K~�I����O����asx��J��XTZ���y�]l�m��,����Q�����