XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(5%fXR�H�����7��F�,R���N7�'R:1����Ѯ �"�DH�>�1�.<p�����
���❘��x#�MU��2��t6Y2]d�Ɣ�������fg�$�CW��a_���
=��x�չg������%g�+��K�!"6����	�"^`VKb�����I:�I9w�7A�P��
�G�T�W�p��r��.�i����g��i�6��~Ϻl����o�yc0 :;V�_�y*��D�<��4�/�H�+���|`�D�f5��#����9� M4xT@I1gy�Mdf�ے�|�w_����3F/7_��z��g�&�Ȋk��}�\�e�*���y���u?i�hl����"9�'�P�]U�m���ޚ������{.9��8�7���@��1�5�°>�X	Ɯ�>�T�;��p�!?QnT~N�ؗ�m��7%�ҡ]T�~��09��N�U�,�G?���VA)��!{\�glIa��#��@�R�H1�j�� .�����%�.vɲ��h���#_ܬJ?�ZS�1#bDm��[yPe}W�d�P���OacJ6=av	KK��Gk��0����4f�v?�=1��`��(�d��:L&��?����2�*��(�Gɓg�>��Hb��SΨݧ�F��%��Rmͧ^S*/3�Υ��
Չ�  ����b���۸�ݔ�Wu��tv��ޕ��5/� ��_>�ܦ
&�Ȕ$h����u��*�:ZvB*��Y�4���!Yqp{h��OXlxVHYEB    fa00    28c0�v~u��lY9;Aj�HdB��/�����~'�産e�ޅ��j����,4y�����W�>4H�UvN����{�/�p���r�r�m�v.5�����HN�"��7-��Y��	+��1`���~�����q�{�	if&��s��lrĀ�֏�N��)�,�"��h"��Z�0V��Ŏ	��Q�9����Ŷ���]J(6��!�g�<S4�WL���nV���`5C�8 �҉���F!zN�M_�� �Kl���_�mp��ѱ����s
m E�X,]wi(�6����j�k�js����`����D ����s�V/��T��T������%��_�1����σutנ�+�4���� ���#�NF��Y�y�`�d7����!��<����'��	/�A���A�Fn(15Y�f�?�}��,3���U9�܆5���%�Qpv�>��؆A�.�M��Z}̘��@a��c52H�U=�}���&@����*���>e*#��fBZ����özr��O�t�Ͻu�F���AX!��H�������y�A`��c����y���vE��:I*M$�����Y)S��쵢p.K(��]�i&2J��S�7RO��hG�|���<��E������(0����x��P�Q�t��9},z��5�P2Z!�	�	&dhw r�\�V� �i�2=fc�e�k�܉4"no��;���VW�h��=���r��=ă?��SX0�,rQ,紸 .��[t�.�+Hm	I7�I���R����^�sJȡXuh1(�P��xq1|لp��d�g�]&�����������8<z�%`�r�:��gog�׶
cb����E�$���2ٰۏm�K�_�5�� YS��߂�'�ski�;��}
̶�0�[_�	 �J�gY��X- X~��p�8�~�^�1���6% �2�mzN��D�+�KU�q��?;踏dQAؔ����]$d���Y�T��8"\� �<�;��@Ƶ��{��Z�?؜��Ś�"k�K�ۮ����]Ù.j9 �����K�����71��N4�÷M4�_78)��f첨��=���R{M?�]Ku����~��T�q���(���KG牚��}fo��_3����X�	@2{��ۢ?�a�o ��<�ө�v >�������c�J��z�}�@.o�Nِ��?/N����x�QпF�!��E����B���4��� |�����6q��M=�ޕun����sge��S�}o��[���1��%?�v�\�B5XrH�:%�>!$&���Or*���^���<�����e�c했����ˬl���w��1$Ojĺ�¡c÷��X��]���;���접���(��?_H2 ��G�dR(jc��W���)n{G�����K��=^����s�w����-j͵�Y	�s��9A�u���j �g5�ҁ(�M��P��~���U�Ӭ߯���l9�KY�d;^���!�!�9�F
�A�妟y���`�R)$d��@���m�
�"�},�0M�/�tS��J:;��hY��ꮰuVpG�a�uk���>h�_ ����g$�1���9��i1���-1��*�<��N����6�/ b,��4_w���ĺ�(�!�%~�U�������N��ז��2&A.����^æ�B��=?�lw�(q������ ���p����<��&�E��E�zզ��]ǫ�-�a��;��U�g�P糲��i��\k��C�]�k�&4��d}�l��=VKG�l|qe�<E�*Z�n�[��d,����lL��C\(7�.jܕ�Pt8����Eh����M>n\��7 ?��o�.t�?	��$�K=oݍ��E�J}E�(��ZĒ�}3QE����ɫy��G+%����:s���l�Q�c�a֫��X\��o���*Zr�Cf�ר1��x�N��]R_����5{�ݙ��F"��<���93�&�n��aD��NK
�ކ������03{�ؚA����$���l�>��Azx�+kƉ�����\��y���#���<�(0T����n&���.�K/{R�J������4l�s	�xXt��j�Gѽ	Ķrs�FiK�o�G�|�?�����Ǫ���!ē�>Z���mIvxb�M9\4��@�8�8ٓ���=���r��pց׉�^�R�\����7BlV�#t�D��е-�x�TA�k�z�N��������c:7Fg�T]S/T�����#ꧠ�N�L�]b�57��{�����q��v�v2��L��>�!���.|�͆Dl����u�x��|>4���ʻtDz%*i��4��E8c�fzR|w�F��y�Չ��al4<����b� ��R�r��	��j���%iYlra&l�a&|��Ǜ��?pwujȢ���Ⱦ���36��8�����3�e���z����"|�*	Q������"V\�3���wO9��_��e�!I4_u� �gң2{���n��)ǡі�S���	�
���S��I��n�v�2�Y�����i�1V=���vY�x>��8T{G���U��@޳��;u{�
����^��H"�	."ˍ�L�[)�/雋�c���K�;�408j|t�mi�	F�N�{��Y��<c����Θ	�X@��iK��Ek�@�{yV�i���J�����<|�����T<��.���U����`V���V�>���xh�oݯ/#Bv֞�a$��l�]��r%�R�k<t;D��4����3��KqU�ژZ3�w4��"X�����y`��m��t��3�k=)��d?n��+�I�L7�ض�Yd��;��X�wA�����*�s��9�EZҿ���ʌ	=����T"?�,�qٕÂԠ�q�!U����F�q����!�XZ!��C��ؙذ��S[!����^��m�`�BSoL�MVx�\"y�IT��5*�����j�	
� �v$�p�P�e27�%�a��X����G�#����܈\$/���M9��TB�2S�6_�ԁ���'c: J$r�T;1�Db;�m��a���!-A�++���h(�GQ����1e?�t�{l�5P0[�_7��-S�ҙ����s��axv�����Z���d�"~��B9E@`f<g��gV�2�.c�~���h�#�HT2b��҇�V@Q�5Zj��:�t}|-���2w��i8�������+{�\T"Y;~���fW=��q@�d�Q*T�@���G����HcCC?Ib9�5$3��(��L�m N���#��>�R4�2��@z���&�3����Ҙnz䖿��ﭫ4�w3Pt���[U,���֝���+"�����m�-&(V\�q�	�"�v�0���߹���/���<�-@_��m�����X�|��1;^\S�$tj��:��S�aՌ�p�y)(�ZX�.�x����Lf�vǚ�zh�1ˍw� ���%�}���Y�g-|WW������i�*�����V/�������d|B�o�Y���p3::J�K��]����C��#ߠ�Jl���YB84w���&�@��?h�A,˓��>��EbshD������I	��0�c���dP��?������Gҙ��t	���2�^��B(s¿�e�+"T�3	}�G��d�s��mЮ�f$�Ug�LV�k�|4�E�T&���iZ���y$���@�pD���Ԏ��;S'c���<�P\�ޮM�,�L.�zm��5a����S��$�C�}���k��+P��-p=�7{�v�c I�I�"�\��>�Jf��N]����P�緸1WCu�wKx�(e-�=�rNo�ٷ�|PJR�8D��U��ƅ��� ��B���f}Z�I��}&���jO��'�܋H�,:DQ��ԫ��\�p12�j� >Gf��5��)"Q8�3�>NNR72Y+����}�ӢD�ش�y���{3*��Y�K���7��0����_�Vo���Z �����%苗;����B���t[:������aF��br�şmb�5��֔qo���#��W�%0�cs��\������c�YI^9�h����� n����:^7�N��"4`@|,�����9U9H�	�%�UV���H��݋'	
�� �r��I�]��ْgH/�n�eY�g��W����VDm��4�$��T�B� ��qV׮t��X�l��C����Ӓ����6&��cZ���P�[�����7��+(�U Ϯ,�l���£����!@�F��x�^cG�����9Է�*L�4.��دg�~�{�t�L���;���.]ȣ5e�������U�(8�:{�91e�jrkN���F�6��A�����ޥ�~̾C��;/V���;<1�I��F� n�}��M��d�	/xl[ZB1m����	�7苨�^�P����Y^_	;{~���
�$��~<zz�S���G�Rw�0�/�i�����ń:$?����1�e�6��K���`�Z��{?�׀�g�Sq��^�!���g�*ԮdO,R�޷=E�[�⛫��6�:���јĮ|��Z�TB�B%)7��@�G�ޗ���s:�f掕���x%8�Զ�x�%ĵ��+�6Zm���N�`:ᓡX��T�P�,���=>^�ݑ�ٕݬG���J"��,]W�����I�Ќ^��9�������_t�E_���eg����Pi��_��$��d��p���ꃝ��[?��tZ]�:|��WZ���>�q]��d�z��ZvK[!�AI�Y��J���xh��d��đl���zp����-��K�֑B;�DV������LUm)�P&'�B��$3�Q>_���5�O����sɳ��h��(�5\�_p�>�$�#��p ��l��8���Ǧ�ml�i lӎ�C9H�㏟V:I%���/�m�0�h��-��N�O~ ������E6}ǒ٣�$�/��7V^*GC*�9�J�敗����P���Z9�{������ǌ��MB�?�P/effzjã6�(o�_�Ǔ���NP�;PF���Z���?4��%�9��Gj��	Lsr.�2lBoF��d�Js"�y�A����Ҧ���l��qۤ��ĥ�����Œ�Sۂyt�njn��׫4WK��9��^Ȧ�x�7v��)��X���?{d���>
	�!{[{��z?��v����è��>�2�֨l����VA�oQ=6�j��.#F-dA����ZN�x��	TŎ��	ր�K�����Ne�9����,+3/t�u�)�Z� �ҺZTއ_��ٱ �?/�P�W��ݍz��׷u�f��M���b�����<�w��CX�wb.�x��I����qbGj#ͨ��<�Ϭг\��}��{*(V�]�����x��������S��W����Py�~Iۖ�5.�(��4�Խ*W'0���N�x�\E9A�ߍIp{1���-l�o���ˬ� >��K�Q7c���`�G�xɞWV�����6�8}n:����I�!�@v�P�R"����hG�Iз��.��յ6PǊ�:��i}�/���	��#S&��
���͔w��G��UK��֕�����W��q�*R�b�߅�^�=��t�mW�����>�`�!u�g&����Y`��g��}�OK�!���>���]�^����`RN$h�C��ߜ��PmH��Ө�V�ҳ Xc��9H�*���͵IO:�-R����o��#`M��s8k���h�V�n�L{���e���|a�8J)����a8�ڰ�/,%s���څ�'t��O�:�߱�ٵ�U�^ܠ��&۳�����cs>˹k0��DMd�3�s����7�3���S�0;��er�E�o��-�d/�P��['o����ys�H����M]3�������Q3�u�t�lo��L�Q)�ȘG�σ��^j�p���\�}Z���䒀j�͑�𙽙��&��D�j�n�������o�-f��0d&�%��}�:��������&��w��	�^�����8�߆�菃&�H\��g��Z�ʫ�,�����w���=��:�8{w�rb��T�ef�7��� ,R�p�+��4��܋֎A+�x+]Z���N�|R� �ê"O���jṡ�������Xd� WP�*�Z���(�<���߮�s�'����#��.@��bؤ�y�F����{��l����L��ﰀX�7���G���I�vt�7�w�7;��1��Ъϲ|�ծ��ﻜ�av�]�^ϫ�N判�����h�
8-�iv�~r]O1-7*R���Y���ui�����Y��QiظtM@��`��ީ��)�e2�Q�e�QŦ&IfQӷR`��Whj0�@w��g��@��~�m�$"���)������΍;-��a�%!�`u�}|Mö�+^D�������M:)��_����p�����vs�v���^|+V J�=��O�e�(;U%�QK:�JM1;��arG�Dbbu�>�&D2�B.��;��8K��\0A��ŒL'{W�q���"��*�uu+γK�4���h�~�c||���#�B��⺥G�b}l���� �'�_Q�����������O�g�2��]d5�oP�N�&�T��\K2;L�*ϖ6���s��W��
Ph�*	X����QP��Fl@�G�5����$`�-Z�$�h�C������i��V�ۼ�RJdF��8Ny&x��C�_[~�ȉ_Ӄ$�#�M���M�z���6ge6L�8X�B�N
�rG��^���_@5ՌM��ܢ���&�I<�J����}��i5��?A�Ѩ��ߋ���,E��{�[�0��	k�8�A�qu�(>��&�����(e��]=a����j � �e�?�[t����"��1�J�B��Ӆˤ4�Uv�m�;#�]=��=�K�=�1���.�S�ND3�a-�����Ū�\�������[A%koE9��\��KiC����ӋJ�B9���r�@S���0]pG��~IF��wiHC��a��NL�N�D[ʵ�E�#%����T�I�2�)f�_�Hv��g��o���I� �D:+[ra��&b��t��
�tt����2���T�)��ۑ�2g��I���^T��8҉�����O��y�oQ��@|ux/�^�"�NU;v�N�80���s��,�aK���$9Q�wvL�>FTG���D��FO����H1�5V��T�P�lU1v�*�}�LbX�< /¢���SNveE�r��s���%��Gw��bü����������3;�������&��"s�j�$M���	\p w�R�^�]�E��}W[R�ɀr�RGxu|#��2@��������U��ğ)sK��rU���m��x֨��m���9؟SAX�#��h��:~���,�<�u��I����@(Ԗ�V'�ޝ�V%�x��1�|k&��{��j7���wP��*_��K �Μ���B��;o ��0=.�hT��TtN��=����>G��Pe5g �Ki ��P�<>ϥ��]����[E\��>��T#.�~^ډ��ךsɲtz稻�̊�n�1r�_���)������[K:�C�)N`m%�Q{�m��+� ��
oP����8~�/���wl��A���ߌ����P�K� �ϸu�����i��lh���2<����qN�/'v�d	�hQ�������i���� �cXQ�����Υ)��`]�Z���pH��?L)��@�^'55M����N)�����vM�19vjg����G�h�����L$�<�&buȽa�|=�t� Yj����+ݗ����q�[��=�K����k������^��-N���ϋ��ܦ]'㭳FO�,wF���L���C�se���"�����C�$�'Z��\r�}�siJc��ݵ�i�l�V@�����8�����F�Σgū�d���bĒ�H�k@Q���ZV����q�����;*e�CJ����à�h�z6(1�ߕȱ:��I�e�0�A�}K{L�0�E"n ˕�&�{�����.D�m�@�Q�'��k�DRڕ�FOA�/1��Ԗ"�uߙ��I2��ڪ-T=J����FX�23ҁ�7[���G��~��*v����J���i�e&A%�ٲeJ�O������Q
��2�����*u��16��n*K]L[R��S;�^�:}��Q�)�n��u���Mj4���%g"������}ä}=DROP��8�p�	?�ڄ�������*o%�{D3�} �\.Q�Ie���NTc�P�1� ���o�<��Il��8��C�K�p��������Q����I��Ա��5�����动��C^����4ｃ�(�n��{�\:�$����4�p!
�
R8c��ů��q����[}��A�E�Ax'��J��M w^�K���p����	�Z����o&�Nb������H�D*�8�8�����wH!nN��g���5���J�!E���0In�|�8z7k��Ħ��oЁ���J�[Ce×�qTWk�90����yt� w�ҟ���)��u/Շm��S��G}�	�!�����э������A�"F���.J�76���R�h��B�Nt0�F��d��X������]n��+Z̽�:=*8����%
c[w�_�Z�P�T�?�rU��,�7�sxF�n�!b���8Gl�!}nAbԎ�����Z �K�t-��C���a��+�ժ-���i�{��h�me����$�;�CN��X���V79�j̓;��]����)��,��Y���u�W`�|�<�9YP�5��0,U���Yr]v��f��R�SQ,?�3��{�@�V/�ۍ�Zu ��̇�%�-mD�L�.�X.�n����~����ELV^x�iYi(>*ˊ��[!1�� p�	�#ko��'��JK��p����+�����*���?��n �d`f�k32BIs�C�	�����3�9p3ob�.<� 䓫X���m�g�6_�jP���Y���?4;�c�}�U�^�}�y(�1I���^߷�޶s�i�e?��,�a�-�}�-j�yR�V(@��R��BN�2<<�Κ�N�8�
_q�?c1j4 �����+�Qx�*M�����p�輜h7�c��L�	N�KR���"{\���v�Vò�̗ߙi��s
����>�.���ST�eq�}{�]��p�?7��è�Oh��EN\EOi�ߡ��$-�:p��i�;>e�tۋ�s�Z �T�pF)^)a��[��R7& ]��)WE�^@�}����(�iOB��x�7V�L/�׊Y��*�����IN���H.��*^���"U(z���]Vx�p|��W�����+0�7� P�+�/��=`z/Uhox��nR�)�%�@���d�� ��^q��O�&l������M'9�u��X=Zа4���%��U��a��nT��>%Ww\
�V�t�E�X)d�xӫ�	�}�������@ڥ��)��0٨�zpb����{䵡�d���F#����"':�F0I~�7�@�nҍ͏�Ι_�_y������o��"F^���������*��
�k6�i��?iɦ+#A�7���fh�̭�B�<��M"G�{�8o�~��T�-�ȧW�)ګ4����S-ULr�����j��[MtNG��ǜw�J�&.�x��t�S���?GN�8�@�V��!M����B�>J����\}!]�*;���;O�`��C����7������t���D�>�j?g�@K&���PTd���/�y����˳��N"��Z���F/�2!��O	�ZD;���3}-���ېU��Pm#z���"K��Lj�*Sk�zi�����?��RĶo��֚�b���SH>�V0�>'��}��U��u���ˑA�kѼ
����Q���	`���s��|���jP��l���Om�\�y�^-���/8+�����*�j��dl���;YL�aLm@Ա����yU�V��]���nJ���8Gpu<�
�9	i�� ��m�A����e�s"cr%c8�7R�,�[x�S�]���ȡg���(]�W^�h}��CM6ŵId�u��TВVʕ+�@��~�A=�-7��\~&u����G�����y��5��o��C��׾L��?��0R�H�x�`(�K���C�����+N�� .�ڥ�%Uw����~rh�k1C��a^Jhc���r�)*,*��[�g����N��^��XlxVHYEB     896     280�{��rt��8�<��G$�'�.?8���!�-���\ns&� V��MS��6_n=y揺+Fx����&z~I�	�\�Oa������&'#�,vjhI]�HZ�i��bBRz��Q�k�>�O���!s5�d]�"�r�
I܀�D"��.���̈́�s"���{Uo7���N��H��?c��98��h��Qn��>�(�6we0x��O�`�R~���n[uz�yC&��%���a�np!�\.z-�Z{�U�k�g:%����(q<X���+���s���8�y�����AO)o��-z��Y��j��C~C�Z%�CL��:|�=�7I�W1'���dS�w�ă���]���g���{/�H��k�B�����X�X�hm+F,0�g�q��b��:�:h���Z�ɳSO��*��o�n�/rh�E.��\�������`7M�2�b�p�x&_D!�@R��b��£xWC$#�ľ�d��ajR@q�ס�ʩm4��hЇj>g��d����U��b�c:?���z$!�ݫ��4��%s	������7�u�B�9=g*AW0JA��`z���(�� �s�V:9�`���Rb�䓦YnL|�A�����NŝV�~��8��g�!����8�