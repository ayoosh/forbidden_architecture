XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z9�8<
1�̊Yl�&�%c��62P��ǌR�+��W�zwA�#G�0��1���H$C��l=q��m�}3�Q�B�_|�j���Dq�;��~��?�|8��q��� f������b{�(/Z0���֐��<�
��
����8��d`����%��o_,?\@Z�.}�
��A���5=���ef����Մ��kL7ħ���^�畷B�I��a	GV��r>j$��~�;����Oѱ|��d�9o~=w�.�v&��8x��LY��9�i���^h�Nish|�fu�=��a��«)�k�q��\-��S�;�5Z�����wm���&$
W�׶�8ۧ�v��N�`�ᬯ���M��S+��q�ۛ���za�	g|n��#� ��G���j�f�����96�����.@��m�i)w�lh�����`�1����C�x��Z"d�E�x�w��<-G��?m��-�p����g���j��^�@^�I�|ǅ���z��ϓv�b�?�h!�Pws��N�c^<� ���N4���Hr�����@/F�N�Ta���(�BآԺR}_Z�:��D�|U�<�fyJ;[,w�?����;t�G`���.����M�L�)�'��iX�>[�u�o�$�f��,��V1��埿�F�~r?��F�^��������x^��w���G��L��n�z��V��R�E*{��?ak�<�]m��R�	㌿̯�����|����V�C~��	$XlxVHYEB    b8a6    1ac0��#_�?������e
�N�ݓ��Z��X���m2d�`���׉Q�&�X<0\�f��:��Q/��+[>�����|r,���6M$���%�����i;b�a|{6��P�W[���3j��5���?���ue^﹧s�5,MQ_T8
�)�I�%(������^�)'焞>���r����J��oo��Y��&�	n����<hk��\�d�닎�*@^Ç���|�	{�P�SW�{(Ӂ�0�����<p񘲊�����p�]P_�!0���	٬���fG��	/)�R�f���^��[�S���z��~����#7��E][[XOE���+'�ٺ�%(�-���`�P�z����:����K�Pb�o6]�����������
���b}�����68P��Q��IV+Cr��1\2��\G�خw�˖7q�s�Q��覩�$o7�?���_��#uhy >;x��r\������ܩd� �6gbbo�g�Fތ�]C�J]1,I8��<ٟ���4_��������t1�����Nm�8�J^�s{�\$(�@PMKIq�c���˾���66<^[�bt_R��<�2�=Wx�[�X���piV~�'U.'ǿ1�J.����d��.���VoS���_gj�����{��*�%*+�٤��%-����{�O�N���Ӳ�//�9���ȘRrZ�D�c7�g��d�9n
�f�$'
��!���*�^��.��Q�侫�!7�%/D@��R#o���/�'�`{����e��q�GH��Ų;�?yCPe\+K�a��D��d�a� ]��X)`Wqױ��@q �;}'b{�㭩`

�g����?a���G�!i��֘D����ե��p�������l��V���$a�<��������s�.�(�`Ugo��;2��l��h4aM�z)d����:�����.biT���(\���l�&�!�N��kJ����z7�<�e4��'�G�D�=%2\_g:. ����m����M��=g�h>(=8�K�z�Q��Ղ��4�L2�2m@�����,��~Κ��6;N:l�*�p�g�%�7��@[9�j]V>Q7O����ե`%���!��٧�˅���9�9Rۓ�0���%L�Կ��<	rNȑ���s�8��2�l\*tt�{�nl�
�|f��@#[�f�����}��b���&�����աԺ�~�ke �$��O�K���/�K���gF;r+�wW��P�2�_
�r��E�� ������&�=X۫��u�gR�����
S�6�.A�� ���װ����4���?�}���O�n��%2
�^��C~3LԞ��l��H��E��A��q@mc��);q��9�˃v݈������O.b>u]�`P� JS�ӆe��ڕ�V{S��~/|wŊ��l�І!��T�:QG�Z=Ӝ����5���`�ݰ�.�[:x�j<����Ѷ�e�u4t���Z7�'��N���0��`Gj�L)�fw�[q�e]���>��w�ѓ6�M�a�4�$~
��P����:%]Hdl �����2wlRE*��u�O��J��(�h�qő�o����ͬ�w�@N7�ĽIc
뤰XAz9���yZy���d� '�-�:!}k�?�vN��gǓ�M�_��GՁ&}�e.:V��Z��	�\�P
�MV�)�:l�zn�齨Z�$׋��[���S=�Zw��1fWS�-u�
dۙ��8˛��9o�w����%x���ȥ��]�t0�q#~���� ڢ�2bCHQ)9�I�_"�Fw��P=� n[=�ٟ���U�Sv����,������\B� �TEiX�I��ѺuW|��>:#��cL��6�Y����v�&�d���Il����}�\,��5 ��2B���$C���e�q���n
6v���#�#�|* ����p���k1��L	�>�K��@͡  3�Y�2dF�L�䬁@�m�o���#�@O_#f���Q|#�_Ȍk#���G5�FTٜ*H���BL� *1.Z�
�T @Qy���~���^|_����g�ȫ�{��M�b�Ǉ��X��2�_d���l:=�cor%h�}e�)��ع}B���_��L����f�EΏ���A�b|S����f=6���w�����k�/>�6=2'�1�pd/:��%]��	v9eQ�K�a�����g�����B���������*%�Ӈ���(9��.�<�A�bŶ��U�C�ѹH�g�X��i��2�fP��]�%:}3�n���/��e$Q��"�;R|
���ٻ�*�U�g�d|�[4���;�ւoص�o�מ��m0ϼ)�u���.Q`lBe�"�R!���ܸ��'ٍ>z�☟ ��Ѷy/B8ʼ��(H����ͳN&�I�������ړ'���噜j4��3����'o9D���=MF��*

AFa�5Zۏ����ڟ�΀b<({�AJ��dQ/��{\ZSY zAK��8i�x�F����Զ�K��"N�B%�|(�&��3Ϭ#� ئ�|�>�\�������_4��#L˺��;E[�&���&GyZ���C��r�9����{hՑ4�z�`��8�+�(XS���Ĳ)~/�����C�Y�i�.$������a/�Ŷ6B���z#	�/��7/wŊř�v�c4�ߚY�j���
���`.EE���2<5����-Û��> +��߬S�Bl�{ 8���{��s�א�C�v�9�pI�.z��$�"k�er�Ձ�Ͽ+!ps�ݸ�dl��g�[0��[z��4�#���ܒ�O���ū����[�����b����'�a�]nU�gi��B$��0)}�����=��[b������qxZ�V��S\c�y.�~T�T��z��~T�jV�}4�4�ȕ�8�;�I5g�X����˧	�q"�'�O�[��J�Ik5�X�	�Ew�����9��N�ϱ��$��c6!��/(Ե!1��9f}�$�gU	M z>���I����[,��AY�As D�w�Rx�J��G��}U^�win�{X]�YI����
NA<^{n���>��0����&��1�l��z�t\Ȧ���#���q ��J#�F��Q��MpN_1��w�<���_�q���cr�7�65�W
�~�n3C��	�FP
H_���C���$!5��߰�
�v��Z&�:�� �ۘ�*H��psC������T�wwB�E�M���̑�]�)ytoW<�b�iyfm��Z�o�v?3���m1A�,�/s��
�������F~bi�q��wk�ַ��ud���e��V����2������X&�_sB�@�9L)�x�(�<�3�Ʊ�u��?Np埗�X���R���v�f�)n"�HwɃ��q���E� 2�+���WPk����^�&T�j�F )�^�T��(���ǝg��K�3y8��A�L9��yX�It�M^K�Qo*L�.=��s�R�e�h�f3��G�0�N.��"�j�elQ8���8$�%� ��q<H��Q�q�
�]P"I�g�I�>�������Q���ѓ�!�൲�6�-@d&[�E��%���<�o	�������z
�zWp1�ň?ze'���v�b���2�����-̹l��⸟պ)i�$�����T�\ �~�X��<:�R�(���tEx�{�#�`M'��Z�|�$G`���@�S&B��ǫM�N��$/5)�]�92��J�6^�D3��Ǩ�ń�"�;Rv��D�y6���`���g��r'(��j)d�x���TT�3�W荭&�B��#����k� wװ��]��e�ѳ��a�u>"'���D�uf#O�f��yN���B����f>�t��D���%��`Dy(��p�b�S�Q.������i��yz�x����W�����yO+���
��\����
��2�T	[%�w;x�U�,� �����Q�˧m�h��T��(�ocQ�K��>��L�8��P�	-�I�0+q�r`��&v�r���H�|�i:YP�?3�G�1��W	=��|p�2kؾO@��ʣa��i��޴}�X�i�D��z���a:� �mDn��n���3"x8P�%�DO$J]	���:��@m���P��+0��_�Зs�(�$��^�y�G�>T��˖�m'�JK,,�@�dMz�-c*%z���(�|X�p�A�x��\ɛS���:���5�F�dFi�
������˾@���i�,���H��M��y�y�j1*[P�����}� U��ׂ��s��d�jn�|T��� /��zI���V�澪�华��a�Av��y��]��f,v�$D8X��SC��vF�r�tl��^D'-2�=�����d��<^�*{	uDv����Qm�b���ñ؈�7�#�E�8�Ts�$���|>������ ����^�b�i��H�E�T��FR���L���D>���*�&,��i�0Q���$�#/(��
��ol�_�2�F���W��p=�jƴ�o+�gi�(3w�"�Uf����0����W0[�(^+��Q����*�,��n(�	��֮�F�PC�сǯ�cd�����t�F2��:��
P$�ē�Д��N1uR�td/77�~l�O�E�P*O�����6���]|-�j���<xW�bU��$�F�����Y��.PDރo�|�0��#������+>�A�$�'
�;n�~/M���X;Ũ�,'U�{�����>􀝭�B�DwV	9a�������e�Ş�~�ڬWi�Spu���k᜝"��ڍ�����%HQ�D�|&�#��>�'�����#�t���ͱ �SJ��l�0�y��'Y�9��;j l�����s�g��'Ek�|�L����7��'r��Ĥ���U�̇�l�n(̰��Qro_L*�b��(�f_Z�t*/��t�%^�}�m���=aR����dŴрI��_��4��<�����Vϥ`g�C���i���
l�؃Ț��]sntH&�8��f���^f�������
M�o���&{Iuۛssq�p�Šj2qLҦ��_�|G�h�_���5'Hh���g���gdu� �3�#�c�0�0浈ϐ�w�o��A)����K�Œn�*-�g�yr8���4=hdm�$��>�CS��Mtĳ 86y_�(a��q���v�A(�s���:�-h Ef����䲩�J��$%��sRQ>N�OVۘ�&,�gAAN�4_Ɓx�cTMm��1��{,��X��!~�)P���kNh�1ϩR�Bċz�%�Cs�;�^�tr�����؊/����������邐m��X?�ZС��H"�$Kޮ�G	bE03x�S[6rFz�\I}q�["߮Y]�O�%�Cp��b?>�ť� G�f���e���W [Z7������)��Us�bl����rt1Yyr���I!	J�?� MO�ԯ�(G��^�<�/��IP�W����)oNy�"�2VL�Wg>�%�f_W�
�P�p��g���Y�-=�}6��c��F?K��=p��1m+��+S�5�"� �@��"6h�HIf�耂#�GwsK��<0c+�%2��6m}�����T2�[��R)��piV�,������Č�M���`y� ��*�ZgU��V~�p+̖E��q�|`]&���F,��F��G`�&� o@'�ߟq�8�rLc`駚��Q��/<ݨ��}䋩6��p�X�[���P�f�d���}wH>��f��.J]�>�mA1ٷ���\3Smv��rP�4ж�0}�qe0���7�p�jXk���DD\)���'i%� 8d�*���FȦ�����iި��-b����hU;�S����! V�����'©H�|�Υ���",��'�Q�Pb휚�6դ˸>�3v�=&t�W�3Fy�Y��Ÿ�0A۠2v��0�@0�)\mQ�r�%��jY[kG,6Y�i��{����љ)����'*����(�jr�_���tYY�v���?'���j�z�b���j����|Z�AK��zMDG����
��ھ2�[�oD��g
�=)����"�l~�
͈���!��v�4W=!
Z�@�j�s��#i�H��M!sO~V��ĝv��2��AW(P�j�u\7�{�������?ݘ���B�z�� ��@����D��4�E�[fz<�-Q�C��P6�[�¯�gP�cA]�J�k1�p�Tq��ߦ�,����B
E�K���a���:�ڷ<�W��7(�J�����+��K#�Gj�bh������=9�o^Z����m4���	�R�������3x�ۙ����Ο�pz�M�$��\,���� ܯ�?]��8:}��_�����W�R�J/윃�=�q�V���P��� KUr��]:_�TV	��0��l����S/:Ԇe��0�?|- $N[&-蟙��Q&D2�oZ�w4�7jm��t��KИ�ڂ2�fɛU����eU�'��q�z��l	�Vy�n���{��6��y���q�S'��eϽf�;�	��Vs��<~
�S;��,r��.�&�'YP��W�KK��ww���s����s�T3U�����(c��F�Q�h#�[zs�A ��.��G�y��@�F�i���V��l�iغs,��=�s��\ǿ�����b�i���2Ռ�i�J��