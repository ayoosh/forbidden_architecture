XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T2���i%��s�=�:&>��#w,�B�<�6�S]iv=���e���UB�A�����$�5���?���xzȓ�����R62R���_�ަ��B����{�Y�8+9���#�z��R��T-�??z��"Ll\��"ssqD&�z̍��NP���9D�N�}#�YEܘ^�Q����셃Z���E�%����#����{�����I��љ����l#��Q���X�;7��{��$��4�U��Z#HĮ;[D���MSbQ�P����u�#)�
Om�_dN��5�y.V�-�\�W����������rv�w��OY�za��ڧ�+F.��y^|*;�!R)(N�����Ik��	����5�&�0���ۊ�ɍc�3u��eS�i��9k��q�����p�"���_0W�B�����|�>2g$ ��K0z��P�k���|�� m��ҹ�7��Q�#[��a��a���o",��~�]�Q��L�"�Bv��|Y4[t.eƤ�=�sF��tN���%���ã/X ^MЍ�M����P���qr�n;_
�w��W)���h����RVC�S�IJ�:���Sÿx�9�0�r�%��/��V$�/�͜�/>S'�C�h�1ϩ�_M/��Ͷ?�1F���o$�Rղ.� ��3t�y,8PJ��8��Qw���]�V��8��������P"_]�t�R�"$ǞVq�_V9�m��blZ�"&�:K�#���.�Dm��g�3�Sy���E�!Tn)�׾m�W-}W'XlxVHYEB    fa00    2d60�m��}e;�.�J6�D�%Wc���4t���$ϱ��U�,� ���ÑG�0�u(]�'N�1/=3Q���?$P���)uN���y�8��b5M����6ɪ�=(���F�O�mJ���+�ɍ��+s��R�95)��?���� 5b��J��=j�2:��iGQ�U`p�u�����2&ij-Gl#��ܚ�6���RV�z�ʹ����"R�%�y�H58Uή*j���.�����ȡX�h���v���AiH?\��І�.�?[~2�$�z�t�.Hm��FHnqsK#S/qԙ�w���xra���D�[L��7󑘉���+�2s�����F�W��o��|V:�8<��i�ب�u��S�b)���!�~̥7����E-�I����=�]��,��zf��05\_@\���vbD��,Z���b��'j32�p+�e�W��3���b��LC`�?�#W��I�S-���u ��50��F14�""(ց��U+rJ�N�����G�#�פ�r�ݣ�-���+��,��- Q�ݬ��
 ݻn�0��D��c�NW=������e9���N�WBV�+s8�Y��l��V�Q��@��E̊Tf	���D��S��qj?^N*>��(�"��o���K�
�,Ze���G�z�:�A��:
~�p�A��[j��gVˡL׶>X�P#�}��bG��)[jJ����#��Z��{��5e�USbT��ď��ZgQ��� }ʗsQJ6�㡯�6��W:0�^���5{���)�sW�SL ����[+��"-f���+32C��5�fT�rc���Xrd��Z�l�,�s�"�\�{���O��Z(K�)����*�9��sn֞�R�L�s��P���p��BF����	^�ݭ�_q=��ܼ�B��7�-_@u&�w�^-�!&�zs�},�:��J�[7j/c���~e|3@�� ̔��$2C�UD�}���*̼cQ�[Wʌ^������[�j[R �_��x)�}.JJ�7�Ɉ���(��E�d��]\�.�����qj��N5�Qh��M�����F��E/D�1��%»��4�T�1���0�9�m^�2<y�AF'Ω��_i�SQ�m 1o�a�*�\�H��<�85pq��"��b���"�H�"�1K��!]�i�\�U�h��p��ġ���T�����z��C%*b�0F���`m��QJ�F_��ظԒ)���[�L� �8
d�7�g����wg�x^����8"��7�p�m}��V���tK��Wg�/
wӞ\vh�qa�zn����h� ����#Q��t��8�V�_���`�xՎ��㋋O��yC��G@�<��B#�|�Mg���u[��5�Ye�߈��u�a6A`��qxk;��K��Ǒ���ަ�)���e �^��d�9�$+�t8M~����1z4� Њ�=�;�r��ԏտP>\H���ƀɑ�(u�`�T�I>w��\̺r|������=�0�b(q�*������֤Ύ��7�6�\=�.>g)�.�-Zm� �zy��JI���o�֋},̏�,i� 3/�lm�J��an��o��3�>]�)q��
�m�!�)�M�>I��rZ��ͮ���HIa�j�Ӧ�����^�5�����<
o�n�\���3/����C
Tb�CP��Y�d�Ʈb&��(��ٷ�o�}�5��7�)�1�2	5�� d���eeA(i��~?��E�V�cR��/N�N\홧�{!�������-c`pk�Q�����:~#�)0��1|$���EK_�u�o�l@@���nww��z��qQO���Zk
�F/�W��ƻ)��т�8�g�D�������]�td>����[�tc��;�`�j�N��b�nư�ǭ���	�
^o�2�k���)d_�����F	��H���y�Zq�?]�v�J�sB���%�I� 0��4�H	a�@E�T��; ���#���8��3[�8��r�,��U�R������P�7���2���%j�O<g��?��7�<����S~ί;����Ub��u|ʡ1�`�c�E����z'׃h�c`���*�9¬h��hp��"C�P+SR�j�mE{���`%��� �T<���G��C�{DKHl��8w'|�3��b��0-x(�ԧa-#��OZӞ*; ;�S3�?ŏ3���)K����7ENuvك3���X���4D�w@��W�����@eq�5%�km���.������w���뛁���`�1�g�V�C3�Q�i�I�]c��P,�O*�l3��e%)M�y����ˊ������e�e`�l�Tn�7�%�6IAcmG�!��Cq�����G��n��+\�L��Y�Z�S�h"^>ː�rQ��Tރe�(�k��GdX�W�I{燉��D,<�V~�`H�Y!���CP�2]fzm�����?����+9X0p7�(�'�����{���t��0�f��}o���W9Z�h'��=�,Pt\�L��S����j!���fƉھ^���z{�A7m�<���Tt��Ix�k.���ֱzh��jS���1����b�x&-ȨN�2�� �Ä���8��V<�zD�&�P��� �E�lL��0}��}�	�����Z�@k���hE�/�S�2�Ro�����Qg��7Z�C�נ
�{/S>ms]��1 �A�<�Ε�f�wj��̺�㈧-�8��������������=�	"N ���M�*�Tq��I<���zL�b�i
}_�4Je��O�>�-%�� )��N�1�v͹���+�r�:4-��I����n��M�r���H�C��&��\B&x��t>�(cb��ҧ)u����-l*��N1�܃�ﱬ��*��㖟���k2+Lv�$o@V �)P���@R��Ygr�6��DE���s�_t�Q� )��!�i���UP����9� �^��_�VjjHe�eX�S���'d����-��A6b��bw�oЃ�B������`�~�%.>�����j�v�Ε�F:	7%�� d����@&��v���W'����x�ɸ�;Jlq����R�[�R��K~*\H�ujn�����������&���:CP�@Os)H�3�Ok
k�`�kG�;�g���c�|�U�EZ�HT�!4V�z��P<`�{������Ȕ+�i����iQׂQ�B�>O��X*#�=-u &	�c������Z��Lf�4��D+(�;=����.`
��y�L��e=+�tt-���Z�)bMO�s2C��Pc'!�*:��G�n�k�l�Yw̩���9�r^�,����8���YؒN�N����U�#Y�4Y�t��u��Z�I�x���>Љ�!W��񝧋�S\��ը@�:Ъ����t��_q8!mqd�`�	�6��%���ue���4'��K�<'�̔"r�8�����ߴN�7��2Q�L[W�'�^�n�j�K\�]��]�+�:{� �v��1�u�핲���R��U��z���0��G���[o�Л��L+�g��:�f�*��yP��	�C+��"��8_ff����6��������V7ľ���K�&C�gc��o@ޯ�Wr���Ãs�m(v5�z�$�}�)F��ƜT= ��ޙxz��:�A�*)��z����O������1;2t��e��+�j��#Qw��3l����S��$DTl
�s�gt��Q�`�8���޻;�{�q��L�7c�u4�0C��TLߵƞϏۀ���"~�N��<a���(7!���v�J�I.������p`%�ykRR���Ĩh�q8�k��4���%��_�*%�C_�R�x�iU�����>�)>�a�G>�嬁쉽�A@�jU��-��gq?:�
�a���J1�-�a��h�d��L�SfNn$(���/�����BL��Kh�+Xy+���]ĮL=:H�l�L����F��W�ZW8��������Rx�++�Vi8���g�x�����W�J�9�=h*r�����_2u:�f�ʉ0�]�5�\IT�
�d����̏;{�N����L����
%Y}��ȃ�!
	$����L��.d�2�����V�;�Ʋz�b&#2��W�-M�e�ncb�G��yөtd���5�V��D��������!�_� �Z봐��6��[ђ�T�stEwhv���"��n����`���n��J,7L�����)?}<LT?�����x��^�68]�5?ٿ��M퍄��A���opqw�_o=-}8d,��������$W�Y�!�MF�z�rD�}����P����1�x������4I���X���t*�S�-/������%���tqu�z;�$����/m��zN�U��~��� !7r	!!b�~�%��>r{!?�J{�7z�
I�g� ��XN�iK7wJ�_�ۓ�%d��*ԴaV����l%1����z���EN�yМEtE�s��7��,t�P��l��P�^��֒i�><�z\�
\�� ��M:���Zn��IU����M�e�h$�"4��U-�]�
����9�Pr�8�>�x����P3m�N���s��_M������k�N	�GF�Z��\��ҁad���
աď_]Czl]U:E;��)7�f�H�K?<�����N�e���
�Z�Nf�uH�v���0�����n��2��2ΰ���?i��w�����# i��v������g�Ѿn�#�
���;��{&bRl�a�f���٤��TG@18>}W|&�.�^�G��[bD��1,�&S�o�X�Ƌ̤J1%?�O��k����o.oS�u-����׸kB��X�&�YoSO�~T΀�x&kR���@���yw���v��6�왍�h5CL�5u(�KbE�6RZ�+����3��1�/_��d�X����<�qi
X�'��0�?q�mp�?�&?�L��c(:8Ģ�4���Q. ���u�$l͑�V]�s
S��5&S!_ܩ�dŔ�<�B�Q��zEP�Rd�}������'��? S�Q���d$(X;?5���~�� %�q]R���l_�b�p2�,��Dt*����*G�_�a�2N�j�H�$XP$#b˫��C|����F��h�s� ��4,��0���:�b�K������	*ז8�����I����uLt�g��1���F��ʗ�%�V�֋��܁��1�$|&�A������#%�&9
���ЄB����=dg�j9,���W|_Ō�D<���T	��6!�C�Oأ��3'��P����y(�I
����\��|]H��n�m��Z�%;�W֘R�qޔS/4o�l�3���J�<���֨r*!/k6Aeyߖ�\�A�-'<�S�=g~�Ul"a�h�6�I�Mh��S�R?����=#�l�ӌ�
"����/;ݣ�'.!�R@Bx��.)e�<��\j-�s�o�tmY�l35r*�sr�h���o��#�/>�ʸ���bY]��92j&1R�������{�$m��#5ڱ�	���/Sy�w�	D�Ǚ��4!>�<u6�7���H���,S�)���|�]�V�J��|��ų���#d��ug���� �85>�������ω֞8�}*}�['{�-�U���?�'&"�BI�����i�@@���i�.t�r^1�ނ^U�H
����+[G>�>s"��q��F��L�_�����Fs��ڋ��|����ET���F�X�&^ա�J����f)%�<QI��]�H��|�G�����J1U
���	�����ģ��\�K���b<�|��rwBm��@��Ж6���4���R��r����,]�0C�<�B�J�nŝ���>�(]�v˲�t_]��] B�)f�K����cj�f��4�8�,��h<��o�Z��I�!;PؗL� jW`�8����H����V�ţ�#�g'{��`�F�@X��!H�Һ���bkS�uB�,N2=��y���<{.1�o�5�Ҏ1ߣ��sP�E\�i��"�?m�ȩs������w�`��l�bp����4\j�}9tq�%f뛖A�.r�e L��|_�-K����`iN�7��\�Y��E�%�,��B���dѨ@�ԛ�פ�N/$K�|�Ċ���aku
�@c���5�r֔3����'��D�Y؟Y��:� �.�
 X���T��/H"��~_��0{}�֢�-��iG�Q�����w��=%��IDi���+��3��������.�Պ��qƴ1�Z��G�x"pb4�5���d�Ŷ����K� �#n�b�#� \�J<�q[�i'�w!��հ[8/��'~�=i�JQm�9X;�d�Ʃ�z���T唈��(�A�bϧ���K�t��E�_F�
�u������?k(��> bf�nAi�,u��C�R����@�)#NKY�>���/h���S��g��7f��,"�Yc{Wˀr`3�t跷M��Y����L�D8�G���a4�4�]6�餚/��EJ)�Yu-���S��Y����~%&���>�;�G|Wj|��n��G���66T�J�/��+��M�H(x��|�G���CקXҜ�t�	J�:�;�ѓ�RJ�ʑy8�O�Wo�gA3ǒ�ԷM�������u���ޟ)��?���9q��w������%�=����p�.hi$���#%'г2��T����P�!��X�����v�ͼt(���X�����y>ZcI�1�賱\ktN��r8�����+��1{�N��p�W�ۖ���^�%a=�U:��6ѕ���BycVAs-�tr*��vF�����6�u���C��U-�,�-q}CipV���<�}����=�^m5�0�)=P�U&����U� .L�;�8mYIt���#**�(=��[ST�L5��L�Q%�;��� �5c�TzE8���dUpL6m��z)�(�ݡ3��U���f ��5$D�˂���M0/�M�y-z��_��:�����P�#�M -8Dx�Q��g;W5n!�َS�p7Y��$��f���3���̶��9��l|�h���O9Z�}*$�r��lb˓�D5�3�p �V�&:��+�?oL��IkiI ��N���(�r�s��O�#����g���Ph��jT��ޜy��K����dM�.�q�������0�o��	oH�Հ��W���T�9l���p�ױ��uZH�ʘ�4�`���͂����P|K}{��"W6��mdA�+r vJ~�5O+�$cW4��.��d�l�:�J��k��Q�:Z��P7��g]�w�)��k���dC5���o��C�a%�/�����B<S��@�� �m��Z�ҝ̑>�b�ދ���AVQ9��\7���Ѵ:T�Ԣ/��	�:W�S���P?יT�U��p�"���/����E�E;�ݐ�n��6�'�q��Bl��mC;v�	��J�5��\f���z-9tH�MH�	������RrBr��L�{(�13��3��#�#�]9&3�YNaэ:�-gq.f���Sج ����Tޯ�Uw>���~t"�FI����r�C�D�M�B���?s�(�K;x+�0�lQ�J#PAs��:������!���pu����������X:�n��1��� �h�Z���yJ,`�
O�oe����K)\� �y"$���h�{ŮG���Z��(E �wn���N���{K�w��[�+ ���j�W�fc3
[t�&�C(�|�[$��~bt3(��؜��8����bN�q����	Id���e��؀R�	�C4�fc���'B ��o&#i�{�<�'E3l���Ć�^%����U���<�Gs
v�9�m�~5�)����������q<�����1�@(04�i��p�>�c!7_��D
�*6ϲ=7����%l���Cj'ȯѝk�c%� ��Gp�6�Oaq�0�0����@ G��q��fmi���o�շ��ס�÷S���6KP��nn&N�E	����!5@�La�K�'���u�<����?y�hh�0,��UJ�5:�F �kz#^�� �yc���V�o2���."�;m�H�J�NU��H�%�SCz�!��X�,��I�=���snه����s�:p[�����?j��/����
�kx-�?��>�oz���_�ꚅr�_9H�s}��ؔD������҉�A���~%ݨ��'��݈\��>6��%,%z[��})Z� �cǵ^7'�DԚ=�~v�����Ҁx�$��&R���<۫����$T�jRb�R���(R]Z�s�O�f�)'j%�I����N׏��I<6
����p���.U� �ė�JA�I����8VHY��EJ�)ٚ*y��0~��R����Q(6��0���r�Q����|�-3u�k����o'O��t�N��AHeG��I�}�m�̚#,=�al(�y �#���/��d&�?�L�Эܗc����q��PA��8]�	�<��_;Xi�,a�5�u�l��z��[e����
n: zP*�2���al<[�Q7�~9�Lxp���$���w]2��<�^@D�R?�l����%��������y��v���#�K/�
|r���w/ٸ�Ӑ紆5�~�}"�+^����3�%���7������<H&n��jN�	�޷�0�(u����]YL��ͻ���X�ֺ���蔛��z��ob�"]�a��beF�c���䅠X_(�� �/!w΅Av�OG�4��^�l
���*V��;�+�.a���͹����@�v�^?�B!�V�ePu��ꬃ�����r���c�4�<&Y{�t�B2���-+�#�RK��Jt3Rʚ�?u�\�v��+�̣?B���xD��u7�N����3S`a�*i�9����yL�I��k����>��#�gJ��u���i��*p2�֯h�0�����Q��X��ƶ=�c.l7����Vj������K�J�U�h�Cf��u���(8�X���E�	c�V��.�<����	����X��zq<��*��U�Vq���D�Z���"�y˛��k6S~���EGa����\Kt�yw��R�����6�{��Ě9����p�xT�"��r�1)��.�>�o�<�sw7�x���x5�עz,Иk�؊5j�t<��a�yH�;�!B��ݳL��,�����=��������$������]�$_?2��\̡�T��&;��Nn���#�T��ܓ�C)�L>���,M��4�d;�� 3�]@�En�Cw(:�#�1�|�����TE�D�u�YC[a�U�����6��Q���ǘ�T�tKg�0�b&��/J_�+��7j�x��ې��c��\�l=���^�u��������jc�t3�3�M��Y�ȣ�ws�K<g_�_=J{��H����2C<ׄlV���Y
�~TB�Yq�?�~~u�bG��q�m5^�_�UK3 Nf����f~6DB�O��b�7>A���+,7V��7�3K����v1��r.q�O�{�fsó��
�^@Y��=�!=j	�ű��������y�q�%�Hv��F��f�V�+�n_���:i6�ު:��%����'ς�J,�8����։$uX�Ed-
�U��ɓ���h�z��T)&���3�\����{gk���������C#v_�'b^��g��v��O�̡x�yi,�md��n���j�ި�t�I�k-k�59c���‧f뭑�(H瘅����Ge$��v?A2/��?g�G�� M8HO�����fz�s�d�޿Wx��~`=�b!%n�ЪE?մY�'a(�^BQY�n��2jA�[�"|��}v���%�0ӰO�cw��qZLp"�Qo ���+?dLc s��i7Q�Q��O��rF�v�#k�e��R&�3�0Ӿ����	�	 n����ƵIFW��ű��C�D�	��C~���(.�8�����b�@�<��[�${���WM�E�e���u�/O��B�Y\ ����ۿӭ�U��-|:��&���{��C���,�u�!ͱ3��R���ۧ���a�߅��хMѻ���L!I(�Y](����7�D��ݕh1�!���ww$�n9�l��j[��i�[R@ta����׌� ;��*b���Z�,a���� r��x�"�U?��B*8���RO	�D;?�� �@0��) �n��I�+.\��Xk-�jS�ly�sڪ��$U��B/����x��!�~�����Efz�AQ2�,ē�ն�d�潺�����.��'�ɨcgS��G�{�z�͸���*
۸A��Gf��3��89G�W���{��ዀ�P/�,��٧2�r�-n�HR�����a4|E�U!kn�eUY��y{�q\9�M�&b�cP����>�熞��)O�l�r0r�ҭ�VY��=sKҭ��=l�x$:������V1vu�ȧ.�G$�M�D�z7
�v�e�W�K�:F�'0�T@�כ���-�5nA5FG���u�gc�d",o�}2Z�'���?� �"	��c�s�|�'�H�K�`��_��4�@�/h?%�gz��qL����/��[��o��$h�߷Z���H��N�A:��(�hL��m|\U]R-Q#�n���! 8c�9P��x��t"�>�n���OTwZ�k_m4$Dz�&K��9��~��d"�9?V���zM܌�t��B�"�^��}/�.��_`�?ǋ07&��t�t�ˍ<�6��Qw���v
�߳�m�;1�$����_˨�}��!�����,�����19_b�,�$���kAO
��`.�q��v���დ�,g`����1$�zW}�T�����a�R������/����'9�LN�~o�uMwW�+�yk���p�����2�n�8\��=�Bzӽ��a�Y�����Ma��3���p쵩oDQ��ŞP��t@m����\P~��H�mԺ�J�P�E=�1�9�r� }�OWi� ch*��(��z�L�N�h��&悐�}�wV���^]u}�V0�9�c5�Ã9�X2����#�x�a�[��miNx�tgE��O	Jj�M�i2�U�-��h�2U�,�(_��{6;�s/���t��k{�"uI�������j���"1 ����JE�wE����H.�;�f)�J]wU4�8wW���|��՚ +g��nn�3���I���X�}[��(8JOe1��7���l�A����Ԍ8�3e����b|����_y�*p���G���}�j]w����Y>'9��U����|�ג����V���t��,��Ch�K��sA�Xt/_��.&���|��W��9Vj
���Uc�(���bYs{>��|���VIfҚF�Jx�rG����@�tS5�mӚ,s==+���e:����GLL��fg̠s
݉B�J�������h�ܶ�_�2Vbc�5E���XlxVHYEB    5914     f20���~c;j\#�c��� ��(k�eǊ�o�+:�7�l:�M⹃OweX`{;X��Bx�ĘWX���<��x2RM82���S�-S?�S��%�,���b�w
<O_���*���fZ2�����1}���)��i��V�g�M�V�
2��}sLܼ;C��-%-Ꮰ�~�)jC$�:��v0���ah^`����o9��rVHc���k-���5� ���n�l�ja�xy3����ӊbAM�I���˜�@�#�w7O���$i�!�|L�C��z�2t��8�A�K�D�pNf\d�A1�3U�Sn�㽐\a/͖�1F`�>���?��0A�k��OP�q���E�^����|�4_�xFa�dZR�V���jax�P
�잵�׹_u��:҂����K{.)SG�OA[�]����D&�St�&^�wb���b�B�@:�1�r�����`� ��c>��mt�ki���T�?�{UD�u����ثveݨ���an�ev�4���Z���\.�� �y��Ż�nN��h%B�z�)1?����̯I��
NTz�Y�� 5���2N{���2����0Ԅmt�j�;�Uy�^��E��\�c���djk���n�'���T�R&�~�N���M�+"LԒ,_��M,��2Y�9��8�#��|�g�I$����?P_���sx�v������	��}8$������W-���"L1Ʌ�Y4j��P�����w�+�5�HG
B"�?},9���䫶��כ����W����IA"M{�W6��d����v��j��	��{��ɛѣ�9�WΚ�-qY��&a�ES`�m͸���v�GF�b�)u?��B�7=d��q�mkuGzVI�;�WS[
�íVר�Ijv�.q���=_���v����qcI�'�u�\��X'qI�U���+�����VL���0�y]�exK�ZC"��ûl�;���ry��� 㶽���u1���P�`��fd��+k�u�lG��UގJiY�A#�����j6a�o��=y�yeL���}�w�U��1:F��Q�;�&�����H�ե��E	��8�H{�8ݾk|F2�L�l5��*�ĉ�p $#��n;�R��ps����r�����21Ҙ{����-M͚�K�S8�q��`-O�O_7�#PZ��}�U����Wn���;IZT����g��x\R�Xp�|`8X
��C�~/8En�h�'[�/e���z-�^�?�+��6���+�;�,��]J���6�;y��[R�=>)��${j���n��z�}
��$�V:)���GZ���G���#�i������3!s�qV���H�#Z���j8<��"�P�vx�c=���f�$jmGX;�ǿ4e��/��p�HDU98��C]g����p�U����g�nԷ7#��&���k`�n|�w�w�ڪo�E�ʷQ�u8˔�?����	m8��+%��m:��}8{څ8D[0]U��0 �%��m��K�A�(P��ц�;]W>h����1)W�=Y��}{$iu~G���K�CR�J?2+o}>�GrOw˽3op'�U��Ġ��X��DUV4�%��lد{M��G�B��7"�D�g�]�0QO-J6}4u���-�,���W��L-�C���@�V� R"؋��Eb�6y�oS��r���|��|��E���_C����U,s���ll�5��� �W�G�vR��L����Zս��m�����]�տ�>77+o��e�s5`H@��='�~M��Y�$�_���8�{\AKoR7;�����I���Z�����רHT-�4B6
��9�sr��u-�X����PRb�����lb~@�k�}ӿ�{��F���o�00�sM�����^�����63��h�& ��J�F-{��V���5_�y��4GX��G����C�X�t�9�aaj%���`|I�s�5���b�c������E'Sl��Y��폃�U�5�@�c��z_^,8��CGS�O�&%/Ea���lf'��/�Y�Y���	�,���ּ�3�+S�g����Ԧ�8Æ������7>"W٧�Q�)�#�q�VfW�?����y=��j	���D�>�4)h+[��Z��HJ��vw��,Bw�3�rgA��ƾ�hX���38?Va���o�W�Z��J:2�^������������3���A��|�^�D?�!��9U��Z�ا!���abf�(�����x8 �a;�d�}�g�U�Z��ܶ���xf(�s�����+Z3��*mx�|�Ygs�w��bN�?����3���d���w������!�L�`����~d\���D8��R�T��^˂����TF�>��o�6��LuK6G���Wy�|qT�c��R+7yi�$Fi��{�gE(7�C���7�ʛp���al�"SZE�[H	�� ����d�X��	f=|�#�E�tc�E��Ր�,�B3�����!��_^�B��3������@8s��?�}j��qt�C��V㱀�W<�5"�����)�B�����I�VZ��g*:�%Q������F�T�v�c�Y��49�/���i�T�1���7���a�a�����q ��t��cQ���>#���֡Z)[�	 ;;���J81r�<߱�=\�^�|T�`�I+�Q�#8WU�7.������p��O�3Q�=,X�����:�X��/���Zt坷V�M�	�q��t�p�:r?A��(�n:W�,+S�8�\�����	�!Ɣ�t\5�m�䡗i!�v��k+y�%��)�ֻZ}���ju���S���8�B`�f�E������09!��E�T�h�vU3;�[ne��;��z����5�.��7:4��je'C4�`��q���C<2�Q�;�|�H�N��֗��v�!s���B��36p���<�ڌ�\ t�a�[x�t@�#
&�ѡ���N41MPl+=�'N���~]c��$��N{��S�X�C�����DC�Ӣ�9�9��^x|X�Q�l|�iW�PEF��Q�ԣ��P�%H6![�,��Z"��E�ҋS��˹�bfl�ƃ���;n�Je��km�'�Rb�Q��k�_�n:��{�0�~ ��L\]��}W�ZyK�����M�_L|�f��$^{�6�荬 �Q�C�؊4T�yxGȪ	��#��zb��H��� u?��``gVz��?��CY�O����C�C�,�>����bZt�8�V��&+$�8��x.��㒺%�t��XKlK��JL�	�+�D�^z5�F,�@���e֖ܡ��.��9����Y���v"�"�.�B��8���u)�Kf���$��&|��ʫ*p7H�F��tqI�R@�o�
�@�d��""����ShŻ8gC{����$�9�{�]ط���EyB�uYf�hd�9y-Mљ��e�!8c��l&;��Զ���P���Vיc����؟υ�f��*��^]��i4H��~$."��<s��q �!9c��M��) �!�ݕY*�e�̥���+�$*8��bx�ς�Z��~��}�	yl�ψ����S�9���w@��E8D��Iy�D�6�I����5�'Jy2���q�4�
���8O3�.T5�Ԏ�J�ܺs��Y�������ɶ�:��{<�ˮ�
qp;�XKw���%[6O������#7�ߒ�x�j��1Z�D����T?
Ѐ��-�?���Oe����U�:�5gn�)"hь.[��Z�z~��/9���:̔QK2Cp!�:�]�^���4:n�׆,m�T�����*2EeW��k#dې��D���r|w�!%����>