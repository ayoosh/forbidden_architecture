XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t���W	�٘� +f|썈s�l�׿�;���'�N4w>���-����B(��C�P<$"a������X�/e�HɁQ����z��Ζ���kD�{?��iAf.���K)�,爀�bGX�=d�9�	X��w���F��2�}�A͆ >w��~k�\���^0Z�Ki���#�?B��kq�o!��N�[��Ff)�
�86�]<X������1��~`����\V���\��:���w0����Xc]o���2)����I|:�!����_1�+c��C��x�tnqO�1��j�\�tS�i�X�K`�aKd�������@�������^�����0��y�����-���0�<�n3{�^�gh��.�������20��ܑ^�e �2��Rk陽��>�S�C*q��_r@�Z�L��e&}�k6���Q����<�E��jd�բo���A�<CX�Z�>�4{3��/<]�T� R����w0�yk1�S������1xMzn�,J��B�[DD���8��h@dg�����c�l>k����s[�����g��D���\f�;���\��\=TׯW����>.RyZ'ϭ�U�G�M9d��Գ���nEi��S����:�$�ORȩ��W䷔�,F8d~ނe_��t<����e E�:�:�=��+�ԏFߟ7��.i�YpVO�H�}�v�N�
,��|�/���i��%�u�Y8��}�lnk�("��5i�z�6���	JJXlxVHYEB    56a7    1290�N�	c��2�ELqy���@��Y��ڨ��NK鹳���S��!I�!$�Ią��^�]��d���4%�A�Y>"�?��r�j�a�г?��4.�u%�R�����=+Ȱ�����M���@�ӶD6t�W�沮k��`�CG�l,����y�ݾ�i"L���:��kMA KC�V��i�җ�vD�*����v���[�}�!5(��Pdn�[�Ee�¶��D$/�������T�?|��T��7��^�B/I��X'l����/ߋj��j�=���@�rH��N�X;9�)%��sDT��u�.4� ]��=K�Rlۋ�7j4i	��8���:��@�*�/�YӑVZ�ց��T�i*�{{*
�����/�|����A��(dIuG�%So��W�dl��S��_]���IC�������D���雪�0J|��ֱ��7��H/b�Tq0����E��W��7)俎�4��K'(�1���Ƶ��a���L�c0�Y��F���R�{ƴ�j���T���Ubս�{9���w�%�ȃ�z���jV�'sQ��k�	�EGgȺX�Uh&�e���ϺѨ�����b̥�r,<��[�h��ŴyKC]�+��p�����s� ����!����h��2����%���0�������Y�ǧ��ـ�d��oW��/�{�	�����a���ܞIaq԰���:p�C#P��I��ihč���,|�9�[��I�E5n��|xRâк"K�-iq�Q�R9�G:r؃*�I(Sձ:E��'���۪�
a������o�:$1Ydv�odtK��G���Y�&䓿'�j�b��p�E��-p�E��*;p�_�Gp�!n��83s�R�<h�cr��v�_��n���[�?b�9�K�2�)o�M>�.�6w�I ���7#�F�;�/���D2 �ۋf�R%�E�}p��
�4h=RK�{<^vq��J;�;�Ǚ��f	����#i��Kzu=�<M��G��%px�^��W��ȕ����(�_4�Q�[��Q�pi�V���^�\_y/��N�ñ�Y��Q,�3��sW����G���L��`@gIVcZQp���4r�~6��^�)�K������p��)�I�b
����ܔ���K�@gK�Z��hL�Ե�q|�&8���m�v�Ȱ	[�a��4<]D�+��m�c�E@��t^5ñ	�9�S�'.�����vA��0��m�'{K����B�Tap�,�D�ȕ��vM�����j��^�ƕ��ڞ��Z�\n��Ý/�~�x�;=m�ԡu�L�u΁Ӱ>
�ɽb���l
N���k�;���Z᩵�@\̩阁�����#:�Â>�ծ����d��{�)�U�L�G^ߋ�K|J���6��8����CJ�BῚ8h���Nn��D�yI���,��XL7�J�
�6\cs�P�͙_#�Xf0��2�����T���°��Y����U�Lf�a^�\���Y&_e�w�`�B����Fj����m�� (��O�A>��LD��*np�@��aԆ�O��d=��>��K翷����(h�������` l6�A�)�?o8-�_H9xEضU�Df	�H<�=�u�P���b�ԎH?٩��
6�P�~M��)Մ���]8T^f����tJ�3����|ӰGz��_%0�}�DY�i�u�
0���VP��vU@� �rTf�D�i�JL�c���iU�+�:g�?��S��
f"�R�Z�n���i�b9��2gg1�N}/�̄��-�|@k�������X>��	��k,�70���b�6B^���GՔ��xW�2��7��9��i���J�D ��3ŢG6Y�ֿhf�?�<�{]>n|~r�Y%�.���(�_tz5�!�*a0�z�Z��ZW&�55xi�*yѾ�l�MJ�9ନaj7m�WF@1���|6�*N�{:}��[]F�q����ǟ�;������j�)lb�b�U�:�]�Y�haC�9�uي�#j�*���mg�rg��-F���)���`��4abF�D�D#�\/A��R1R?�DV	��3=9j$h�C������*jbD�:�[���O[����ŀ")�w�i��]δh��g@�-�w�>���E[͔y.Z�v�|�"���ۏ�)�ґUYZ��1<�]�������@E$������B-�&�r�\7������k}oAWYA R�?�#�\��GYB�,`�z�2�u1HzS�"~�`8B��̯�Ln��7�·��	�`��6��=io�Ԝ+��IE���^J Sf`yn�!�z�9����b���+q��2����L=�q���D�׿�!M�����קYB!��Q-k�p�W�9e��Mj�|��a���숾>�O�k�ɓC�I��Dr�1U6�F�S��in9� |�>����"C%����P����U�	tHb:E`@��Bi1qXВs䫪U�̥1*�T{ٻ$�j�N[��>��h�y?ٶUE�6�������^��?>.�2��;��7��d)&&ҀƤJ훫QiKq�E'Y���ە�i����	�2��4u�հ6��~H������p�^D�u*dH�����X��#݅Sl8/�� �C��Dq�*�9��1�5 4ӕ��Q_���4'�Q<	y���������,�,�9�8Y�}\�p&�|��T�>�s/��Æ��l �#�=k]���(�F��w�}����BԐ�g�� ?Aό�t���V��@+9�BV���<�<=�N��[��	L\��.M�x�c�ٍOL�VE�EYbp��:�i�C�4Z�1�
s^'n+��c���;�6~�E?ʴ�m�W��B��ǧ�W�YN8l�H�C�סnj�8aB��W˸��U�!�~+"o�5-����3k���4������x/��E��-D�g6Ũ\�;��{i���+X�o��I=��0���5��(��d[���}��*�3��2P@\w�U5�.Tc��*`�����dL���sEP� ����
�@k�w	?|�ݜ���ǃ�����}Q�[��OkH���Ԫ�d	����)���<���=�@�׏�}O��k���.�m�����?���'�)��(1�3�W��>���4ά+�� ��#V0`�r��cJl��I8às�%�~D�j�x^rvA���\�0�XHo�����A�c�H������A!�uj��=����h2	5�_hMu���A&6�5t6-�N��4�Ku�ٺ0��m����)׭��B���Pv3�B�4ʛ'�����S�S�k����M{��\5��� �U�i���yc_���5:t�_�h]���z����WknC��v^�d�3>�?��&���b��5�ϫ
�sKCG����؄���"Q�-��ě��r�RdP��^��N�j+W��~�!y#j>�!Rĺէ�(U�z�-�\����J�rݤ��\�>((0}�f�?Qp�L��L45��dP�c|3�C��	�͞� Y'����ǲH�k�O������8g�>(���]׾)�Ϫ}U�{>�[�9E�U�3R�#�j�tUyPqZ�J@�6ED�c�D�D�k_d��>o%�{<[�L��_�W�=��䘬���Ǟ�
��Xbk9��	�,�k,/YOS羅��bA��K.�"��5��|7���Xl<�������g!�х �M,,�X0����Z�3��x[�2ws!�PǍ��Rk�}l�[ �
�[��U�s�G�.�ɽ�ڔ�3�Z�Yq���?����TXz����������s�U��[�c�3q�3��qz�x�aɨ�lKQIy����p>��`uA��+�4a�������H�&�pI�i*V��T�F.�����F�ۓVU��7d��lG,I��T�A�~��m�sڏ��S��x���_�,�Ļ�6~ڲ�1�9��'��lV[�/�`�wT[�-��k�Ѯ���f���>W���޶Y��Q 6,	a�/�? �쬧����F~J6\Ug+� �o�:����$Sũ��FG���%�3Đ����A@*>�0��B+� ���b��������,��)��ΥPd���9���Y��zRB�+!�2��{��o���#�<��h�ٝ����O��c�&,��4Wj���D4��٠,�,W�"�Oy�e���!���������m�۬C�XK"�l��d�y�Us#<k�u:�b��
�#��e��9�(Y�uN�]ܗeO"����Y�v��� F��n(X������ƥb��Z�W/�����ެjS���~���͌��r�Wސ[���_��Cc�[M���ΩU_b%�ߥ��n�D���5d��:a=q��d3��?�	Qf��@
Ĝ895a�D~�k�ύJ^rE�}��A�N�9�׌��+Y�$�qک ˓�k�i��	��{�1F�JL�%ȉ})Hn��~2y��((���0�-�G��+Bc���V�ӫ*���`.�@ɒ����u��E��lh �[s�bm�x����U��}�fb�=�g7�u�h�+���aM+E�1 ��F"��SE���Y��#�@�]3##�Q��պ�k�m^A3�G�wy;�)7n�}��5����]���������fm�a����ӰN���6��o[�\	j�n�o^Β*��>��#{�xx�����}�5�#�W���4����f��fJ̉N����Z�&�]