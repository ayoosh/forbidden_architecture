XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]#��n�2o�lWdgG��j[k=���b���Xd���;I�*b��3��o�X�0���`
��G52��.�U��<�����P	n��	�\+��k*"M���	�DV�B�g��5bXHޱE8�l)o�HQ:G�{b[κ�0U�1e�=\�;�	���ǭ�A�gE�ۻu�d��לt��]߂_���3��.\W��B�����&��r�ͣ��p{�yj�UC▓�Aǻ�s&�9�
�'!Hڀ#��P��1���b���!J͚Ͳ�h��td?�{�[�yB8�r��Z7��4�0Z5�\�+J�E������m�m6��ڸ�r)!B�*���������yvB�CF��2o�<ྈdH��I�j�"�$1GH$�ۀ�����l6��ˁ�ۊgU�����L��D�Wַ�:eO�d,O�Oy�Č��+u�R��Xܒ*Wc�F �w�5:E�h
q&�t%�`(�n�����ZA�T�=	������$1.�������Z�|Y�d�����N���Jl�ҋ:���`))"W�_����L��\�{X�r�;+9��c��3�ѐ�<�|{��P�E��_X����u���{%5$7|WG. ����j��ϣZ�� ��kbv�Yx"z-�?��*_�F��5��.�Bj�>�@պ�-�as��%N�56�Ι8V]�*�~_ѕݵ��,�&�p�d��^(�u�(@4V��O���v�h�����/	�'�+\{k=)�J���	Xu&ڪ��HXlxVHYEB    fa00    2030˘D�he|��[a�=P��M;](�7H�e����i��vT4���nX��إ����0��"�yy���z'�;��#G;R�'��o���= ���%U?�n�(��O�DD����sYq�[������"�Q%isĖ�P�y�t��`���A��>��pž�Q�W9�#�-w�Wf�O��)T�N-O���E��n<಺��ON#�V���%E�
����@�,�W�e�R�m6�%ͣI�J[�LH������v]�X|u��"�kA�<��62V�Ʈ��3~F�����~��Ƀ���s9S�=�r�����iR�� N�� ����x�2f��j�MRhF��c�N�8 ��h��0���Q��-Џ����Ȝ=V�v��(ޢ^��-���{�+����.�����,Ӟ]}�L%�1��n�0r�vu�}f�/`֟U�t�ޓ�p�V ㍶��
���̬k`�S{a�M{7v�{�vn	�A�'����9{$�-�:^��IA��rB�"�ykQ��k��Ube����ˋ���(���c�h[�v�#X.Ty�YPmH�ĨH���B?ܫ�2�b��ü�[u�@���C28�+t�_�w��y*sQĹ��t5ܲ�"i�Eָ@��*�[���e��	9����S��?�Z�!�6�;�ˊ%����
�-�K]���G�ꐊ����$�u��^6Z��olwu��یr�s2%,�ꝯJ
�N�d�.u�n��A�/��CO�>3������Q�ؚp��	lz�~R�9������}�{^)W�&uK�Cb��ȩ�@A�$�}�\ҡ!J�\���)AmQh*2e�^����[ M�� O�o5	�в����=~G"�m�itZA��q�-k��8�Q��S Q\S��n߱�[�PWMM��xt��hϥUcTb��:��cUG����U�P���e��	���y�ǜ^��FZ��Z�i���<������MY(|��P�yE1�Eb�i�l�w����[8��e��$��͘��ϝ���5A������?��v~B�m���p���պ{�����!K_��;*���9��P�t�𯀳�@��Z��!�#������P���w�iBCD4k{{�p�=���U C��`����뜿^�=�.(��P4A'iuC�
v�fBh}��ݝ�^Lb��G�ҋX#�;�m�y�>3��Ѻ�`˶��D>9&��E��i�y���>�8Z^=��Ɣғ���W�A���
�'� ��Lpg��\�%S��������,T����.iG���v$v�!ar���mfqCZ3�����2�E׊��9��Zʒ~L�ԡ}�����/$���z���z�³���j0�]׼ns���s�p�1$�׽y��5�S�aF�4&LF��������OP;������Y��H�����ܬ����
�B�`]dA�?��-j+3�ݬ)I^V�T��wY��	=\o_��@��5�k�� ���ׯq�Ӵ~�uh��Ґ5��������y�|��H�A]��7��X4X��m��xOoU�PUR���a����A�Cc�'-Ni�-e-+s/ "U�/31��B=��"��nA4g�.>d˷�1��R����
Bb��t#���;M��tcpJ>���q�"#��&� ��3���g+��`�2<�������!o��nmn��c����>���J=�.��5��O�a�]��՝G,Q�A�G��e��e �����	�횵�.��	~�q�ý�낗�
�s�$�&��2c$9��W�¬"m��d[���E˕ZqU���K����2��p�[F�l{k(4�
�(��(��+�jn�#��'�'������\.Q3��S���7��(��1;�m���*��ߢ�*��u��2����H������CwR i���v��"<�̸����h�i�XH �)j��@G���8
8�y|��4�߶�'�����e��<���WЦ�G�S�Mo2{��eQ3��A��Ы1�U���ʈYHgf�eM�/�Ս���Q2�yd���2 1z��TJþ��-=Q S!Ś��΅M-Y�,)@ʋ��:��_����#�����|�*tI:���(��%[��5�=���a���Ժ� Qc\&Ә�j�nE�G]���S��ê ��M=���1�?v0��+.���<�xHp>���$|d���+*1��Ȟmj�������x���:��6�e-b>c�2¿�V�������  k�q��j�� ��M����;�!�C[���K��+�\8F�pr���±VniH;h�8qΖc137�s�	�{�=�)��������1lٱ�����)A�tCHù+�D�`�vv��{��"�Q��Uπ+5�qI��R��A�:�Y�3����X�e�y������b�ɿ"~�R0�2�a�����b9B\n��P|���3p��ݣ��t�L�?��X�d�P�����ꎥ�щoz�ȸ��x�z�b�t�+O1fjh�r��SP�rW}p�&�PC˙9;1�q�d�H��>w���u�� (�����R$�E���X_�m�ɷ���T~�H��*R��,B�X��[��; Y�}����p*
R�ן�\u�?e�`����y{\�ۻ��� �%�}9p1�z�/b�y>)��y#����	l%��I���8���e�q':�F��n�i�|%sW a�w�J��SY:�U��Q`ѓ�Z�CQ��س@kDTp�0S��F���`��9]x������T�����Pby������-`ױ3H�1���j>^:%�%�]��[����=Mt�q��3�VǆczZ�XF��xxŻ�&ՠTV���W��;>k׌	��/� ���+t&ߛ�A�a��'�~n8�8Uy,����-��YU�;�_O���=�G��Ow�¾ʋ}���.aB��{�B>B�]�E.���;k?׆�n����9L�P:�������}�����:9H瞅�$$_>7�ѩ0([x�g�� ��Y�����/���ر0���U�|שf�t�	�w���I/�͇x���CϮ��K������hxE�|
'2��4�C� ?���@�,��Hѻhց�Q� ��I�� � g߹B)�Aۜ��NVC�ƫ�
{ʧaS���x�h3�y��C�[��!"FT5���׬�Ib���.�o�a��f`�G�U`�*\0�J�͜~.x"�˔⻴�d�6#\�]D<~؛�h?{O�B.M-~zȞZ��%�n�)�&�����p�c/�}���π�,���eTu�v,���g��J"ܫJ� �T�tS�+U�0�������7�Q�7�Υ�v-N#5r�8�m�~DT��� �V�.:~�NA��?�B0����9q['t��y�(�SuB� ��ط��[L��	?
m{>�;F���h���7|Y�	4�q[лuy�zmh��Iw5;�K�ww����Kq�'��J�8~Ei���"y��W�.~��U	E]%V[�V�a8�o��h�fd����3�����릜6���?� ���;\��C!V�~�T璠dD5p�A�������b�g">R/wI�q�8jV�7�� �iz�X��+�H�qe#;��I���C��O�6�~�����E���j�x��#<�c1	�'����Ag�%�d�v��+���lmY�e�"�8� Ө��t�os�2�Y�*�~�Ѵ5"�^2�/�����;%�CW����а\�Vӷ�����Ko�*e�܍Pd�o�=�(�_KB-]���j$��ϩhf)ݪ�g���8�ڝ��=2�x��9-��	<�h�s��~r�{��Sn�pd}���Z�kp�����V�Nl�5�V���^��2Fw��7l)��8nO'"�:�+�F�I&`�V8�7,��8�ry�����@O?������y\�#*L��'&�Lrs$>
�������O3M,A�����n4��S��Q/�/ru� ��TP�s�b��;>,�c3�:�<�Ӫ�6��M�v���zh�wd�Ӏ]zZ�d�57�t�X�s��i�*n�A�k��Ζ�G��d�m����А�yBvq'�Ժ�In0�Dt��9-��59�S��}�V��:b�Ӱ?��rp)�������R/9�ψ6�>R;0�����N	h������:���$O��YRl�#5fF}x��2�Se^��W��/����h,A}�kJ��+ǁ�je�sW�%�WZ�����,��]<I~w	�7���\��r m�]ܗŬO�7E����i\ k~��(��zr8
���i5\Jw�ޟׯ1+�*G����[��U�o�S>�й��Iw�\B��2)���A�@,$^���{g���}PB!��>�X����j����g�U<(��B#�o*��bG�.^hXCT>��@��ZJ�,'�5���C���(#[v4Ҷ�復9y�6_�.V�f}�q���Y��a�4Et���(E�'�H�ܹ�ߜ��U�Sk0�źeR/ ��k#�JM�l~�]Z"8eF� �P�fi��E�{����W`�Q�@���
�����/z8��l5>�U���8�%ul
Z�`��'Md~l4�"d����ΣE9��}��C�ʴ�p$��g/r�F@ر���� K��?�י�Y�D�03Eߏd��������s�R�x�T?��G��8	��_Vع+�OlD2*�i7�^0�#�!Pq��_�w<��5-�ϐ��F�DMT~?����k��h!�@��#����&}���dZ��Y�t��6�Z4㑉*��e2W,���ӓ��V�t!�E��ī^s�vw�������F� @��k�P:���o�aSb�Y�*���<qG��Ut�:Pv[����$���m��x��.���[a����d=�����3t��Ik�$����5�%ѧ^7Z�^h��ں9�I�qKz׼<��@!MP��9��m�$(�m�SP��A�b��MJ����b�|�X��#3q+?��.�{*��-�Cڟ�蟜e�C�Ӌ+����5����HW3��2������Zl�D@3`+�a� s��+K�}1^�G%�y}R��o��^���V�Z�Y�ٛ�z U<t�|���Z�4J�"l)����k �u9��oH�qq�+�=$9�:�a@q4���R��3�>�׉�'��xR��@�oQ>��=���1�	��wCT$[kP�����Ww� NFI�8��w�&�</�֒7÷.�+,#��q
�78О�����[%�QjY��F�:�G%�
 nX����tQ�%e��� �&pw���q)p+�>q�g�b�g]���K沤T	�f9�� �,ȊW&R��WG��\��G|g�M�>�f/�2x�ygЛ��pC��!�L`��²�݊w�.�B.�b���[S|W�,9�y7 ����N��ҵ
y�6���Ӗ��-@��cn��@\m�IN;�A�'�w��E���R$��疋�}z�4��F��K�_�LP`��gO�0�ll��=��?˼�����Ga�>%�!��`��O� �P,�mg��W��L���)� ��m��춌b�ݧ�]h�f0U��y����*�������or���v�a`���̙�s��i�P��<���K/�/��<˳l�ӡ�"�A	8�>�>IsJƟ�ˏ��<WB�l�J.4��J3���?�.�;r��]�gg1:�N���n@�M�q%&�k�����_-��?��g����h���S�Ϯ�"F��!=̉�5h$��<��a�O�j� ��R��Qz�!�ed;�ĀN��ҙf�tS�2�@�7�/����h�4RW�hGR�v���k���Q�-�\���-�	>� ��'�+�'�Ɏ��K�v���c�*��^v��P����A�ҁ4��&&�8:�R��ũ nA
�I�ߠ�۴oU]�Rtggw=�����[��iS9i�O���k憆ۯMdOC�y��x���GX6紨UY�T^E�?	O�f�ϰ%1_Ph�5PΧ��F������!�e����8�{�^���*X��M���m��~ąԈ0�G��F�q�V���?t'�U.���?o���{���ވ��_�W���|=֎��J<~�cBQ����$VGy+;#x���l�xE
m?Eө�{���Y�q�X����m�/�
|���7ߊ@_\��@r�,��|�aaI�g
ͽ\���Lo�1����vz69`�;�����֔�J�L�'��󶫜 ?��8`�P^w���*�������1@}�͉���~��i%AD�ӷ�2\�e5���`���*|������p��8�3�/�&��K$�#�M�H Z�A��@0�=GQ/?�Z֑�O�p\C��c]����: ɸ�x�$��c�S�Κ�x���+�����=�1����BE��(k�W04ҩ� ˨����'�v��#��^�ݦv0�N���6�daBA�-����[0�ʼw,�>V�)Ն�ơ��Qq���G����NQd�׊ε#��t�]]VL-�M����x��P���\���0�~;r�8���Y�%~v��P^���I�t���euA��u��cC�y��ݑ�����j�\{�'R����&�'3ܵV�=�)��DO�D�:�e%�0�ř/�x
�6+��b7895����Ag�h�Y{�j�]	���#]bY!&��g�+�jF:�?s��#údÅ?���	�!�^�'=�<�ebE��J�f% ��l��,��1K��uy��$B�\�u��������`'�}υ ��Q<�8)o�N[����?��oѭT�T����q7��Ƿ�cG�p{'���*�p��C����I^����B���b(� q�NC`�,�:s:SR@ �b}������4`5��g$z9"g��Ӿ��w��;d�SS�J�ڸz���0�ꅘ꿍 ���2��$���ش��>v�zF�=�@A�sÜ;f�	$hY�	�N,&��AD��Սғ���Qn�J����4��nCfO�wN����9�t�Ă��<��@,\K������/��������yܙׁ�C�{[���8�=�m	1���/��E��g{N ��h�+r#&���B6��g�pH�Bּꙣ�Q��[�0�>Jj�[h��
9D�'13q���竌� �gZF�y��$����;�[�b&Ɛ����!U-͞{�ΰF�G ��ol���G�V߉k)un��k���6�{��OW�.4Y�;h
�R���Y�x@/�G��G��:�h�x��[}���ԛ���Ut�'����rY�;���Y/�n��c=���wّr	kh��k�(�Y5��=�]�	O�5���:�����/���P�p���n��l�s }�8`��x�bS��3�7$�R	t����w@�a$3E����6κ`�}L�w�.B�e�+�ĦD�/l�k�+��g�� �����:���h|�a��[\-���������6���5a �
G�B���Hv��S:b�&����b��I��h� �8�m�,��U����
���h(�ħ��(vp)
-��<U��涞���?ʅ�rl��AEU5�L�=N����l�x�~��WE�nW��aL��K�H�?p���.h��;0��4U��5���Ԛ�L��So��R�&*�p]��	�9}X@�|}X�}&Y�XД���<Wb���z��a,���j���Z�����ζ/��m#�_" )kN���5��5��(�Mn!TAQ�ܮ.�7:�;�(�������~Y
`�r��V��&累�x��=X��;�H'm*����7���7P�/njR��D���F����q�#d�O�FŖ��Li�M��U�&���ߎ�E�Y���jB��ƽԑ��ϕ�^�ў�S.��z���sr�9v�;�l�R<$ �
GGc�QCK�"U,���	E�t-���v_6�[��ڋ;�{�m@�%�}��˝����L���BJ�xj�ձ1���n� ���yF�l��8�N��0�����ߌ�WBÑ[���V�֖5��G&VfeH�1�$?���U�����:�1�A��5S�7)(��oT��%n�V�r��8�������Dٚ��=(�SXģW
3�zb�|�}�$�����2M�&,XlxVHYEB    9635     d80-o���*Ln����
��!��hQ���b���W%��x�U�"$#�l8E;�)�����Rm%�V�.��l��e�Ɍ�/ >gN\a�P�\�S�.���)/W��}�՝3+�ɿ����HRH�!XSX��c*9��n 1�>o<B9��ճ�FLR$�4]����Ě}N�RI.��@�~����U��QFτZ�KHFy�^p��WI4��m�*�!u�՗������F�by����)e� �F�߫(VD�I๼�DX5��WB��T��5��u3b�(�ՀĆ�=O*5�M<��<��6�-K�	����3���M5T���;g�Eو������/_Aw���H��n��v�V��	bғBw�����tƀMO��t�o�w�)U��N[�V��N��{t��tJ]+�F�+��F�lM`�O�G�
�~�,��ڈ��_�'�#f�9
U�}�@2�<[�N�_�.�L���.�TŌ���=;#8��p�����@ܔ�A75�01Z�I/0*4�F7!�%�|6�=�����������U��|���I>iSai�׃���Ʒ�S�D�Q@�CtX��0��c�3`9˫�xy���Kr��o
n}�v4Hk�w��i���>*���9g����ǆ�e�pWl�!
JdDe�����Y�ao���x��p��
�^K
R�x���lP���p�u����]&V��������Wמּ�9������"K	��XQ?t��q��i��*��M/b��(�0;|���w������1e�����}���)<<�:ⱙNb$c��:b����DS�J��FhΈEZ�s[#�+ �P���W�~OL�@��;T��pm�,[L>�k�o{M�0�ݾh��n/T� �hz7��l���q~�=�x����@���e=ͧ���rr2;����G�G[��٧�����U^�#�.MW�:�P ���ֽ�����@���0<ڿ�3uɟ������%�m��T�^iS q҃;.� ����K�[����+�X��J�`y.L�	�1����*��9_����J�f�̩}�6U2bY�v�gQ�mR���Z>4�|�m��ϩN��9���d֑#X��ccub${Z���P"i�dX�L���e��Lz޳��خf�n(��I���v�S6�t����+�nW���@KKQF8��� ��/u��:y�6��&/����`�{�q~8>�4�Il���������V�pm��-�l�e*���ގ=^�k'��vm�E����:��d�X��n�i�RA��zE\w�S>T����rc�PbҵG��Z��� ���Bau��(&���om	�$,Xi�.7����?l�P^���H��y5��`�#�����_P}$h���J۠^c(|�o$/�&�����o��Z���Ǉ\��I�%9���s&�׷|� SFT�F�}N��>���G^QR(6�<�1������"R�:�".��_�%-����ۓq���1za�@��ɜ�=ѣ��P�V^��C�h����w�D��Бl	�k+8	�bR�������t� �:�mtj�g�9UG���0��X(=�*~(�`{)q�P�3��;�/�ښ�o�ܯ�ݠ5���x���q)��'���q�Z��%�ڗ@�i'�*�����M���ܑ����#��,�&\�?�4쀕�ɂ
�� �*�����'�K&(_8�H���f��g�id+;Qf��m���u��6�m��SXo(v��vkE�n�����@�o���uR;��f�ߒ���,�M�����) ��g_�h����,�U<�3��0���:���+(�g���:��U)U�NlW���S�烽#lwlϪ�+W��f�Tqލ�����i�i!c�f��sN��#	�[�u�JG�hh���;���-�~���W*��C͎e�Y�*�ִ���#���a?َ�S\L����E�\KI�Z��j^ɓW#ӊ�Í�P|7r"z��:k�S8G���(��W}�L2����n6D�ۂ��Q�|�Ů	@4Sb��).~+�����(�lv�|��dci�g��%>��ni�BZ5jQ�4�>�Ƴm?�MFы �6�/I��U��;��{.2�[s�-T���D���[�]�&����e�K��zl̖�}KQ]C˄�<	F�tj����E車
��	ˎ��WΦfI��R?�*jFH�>�G@��1T�&��B-T:��4؆��^�m3���><[&�t�8�|�䚖������lΜ������%���.�A��[�Y�u\��SGVQ��Q��wY��<S*38��M�Bt��C� ~,./��R��Y��3�������3]Õ��~�C���=�A\K,���qER,�$�<H>h� ��e�+tk�,����'�nAPpMDyr������EL�ʄF�؈d}Av^Km�#kF<QA��w�+6MC��Yy�,&-pޑ���Z$�T����1ۑ�7G���=͹{�{�����d`����ˎGg�}��j�T�T�"�y�6F�F\t$�r�2#,dQM>��W�d�'bCk����M�u�>��d4�l��=c�i��ɲ�3W��3	:��Ve���������J�@�u�ق4ç�._u���b٥ӟ%�w���s��N���A�u��M�{T��|�h_��z��t�f�M]:�[��{�N�(@.��EB-t���ae%�2{n���Ѐ��?�((�����h-��+q&O�d�=3��@�OK�5cX��pw~oa5o�igQ\]F\H�U&XPԈ�[F@<2T$'b�p)�r ��2h�(xj��AQ  1
L�1�r�����h;y��������NBO���bWznxF!��i�
���O �� U�ߋ�d�'�N�r�De#�]p��=��:_�WJi�{l;��#0��o��⡻�x����N��%�H�t�`�>�Q�P��G-��o�	�=lB�l]"�ͷ��0C���F6�cʌ�_��}w�/�=S�'3��f�7��	�s�N5�P�
\ �[�ΤGL�����e
Y&��я��� �[�6�[f!^�x6�ƨB|���Ԃ�e�������q���A&�Ӯ��Wjp3Z�,���q�I�0�t��I�^r��;�hh�Ca�y�LD����A@PCU���?V�3�s[�Λ�A�h7��w�^�tt\	{�3��`jY��_I��m�M��Z�s*��p,�c��L�X3D#�x%�Z!�7��-�
}	C/��� �1�x�)���'�O�m(Rd��*��%�H�|~J�v`����=�wTX�4���'B��Wȱ�t�_��tE�6R^�Y�h��=�&muo�0p�r��K��A��OenBD�C�w���=Z���Ӻ0�ղ�KIAA���Y����N<f��C�G��s��61