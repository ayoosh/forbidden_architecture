XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����|���~z��=����	w��������5���Y��еy�X-���MS5>>�l�K������&w������1��h{�]UBTn�8xb��'�&>��k������'Xڬ8��[Sph�iA�G�����*Mş����o����ʟ��q3-�� f

����6"6�;(>#@��i+I����At�u+��x[oW��E���;�"� S���,s�\`/�������P�CT��w����=���b��6^Q��,5��2��>g��&���J�Yt����o�����>z���WQwsG@'�;���L<tE72r���Gt�y�q��
{��/=�n2KƑ�ȷ���J|�d�
I ;�ZDSk���%�~��OTt��yޮ�g�Ty�]�r���/��E�IE��)8L
�_�mf-���k��!���l�N�������\��!��9E_yF؟YH�W���?��=��j��D�0lّ�>��:��;r����h��f�2<�:]������$�/�����A�O�Ww��Zf�ԋD;�Ɲ��YP-B�����������)TۑWʢ�����d�6d�ߴh���}�x�Zz���������Ȣ�2��!a��z�o��&�ưxb�X�+x&���m�Z�U�~��n�$��Iv������z���`"UPg���oSG0��8�m�]]��x虌>^'q��\DS|E�R��@r��LJ�����H�]�YXlxVHYEB    fa00    1fd0Omݾ�վ�[��Q�o.��0��œ���Wg�^R]��@��KQ������]��2XCq� xG�I�#�\��4p�\#�.e���"ϔ���R<�cV��P����Q�OĔ���*v���/9@b)i3:�C*ag8���1\2����}k?`�[C�8`����>��V,g�=[�� ��<aJ�<j�M���o�s���j�ŁO!�ۅ� ��B���P3/)U��RP��*l�>p{˫cN��G�: Πe�<�#Ԥ�ӌ���,�L�?I9� Pzޡ-�e���ӻf�uQ��RA��7�^���dD1hmb`)n��	�7�1G��!�_V`��_�s�$Kr:��mi�1�F�K̆3/P|Ei���l�������+ு��>9�%^�c��^��a�Ua]�~��Si��2�b��2�#���&mg��&>��,��*.6<��;�$��7"��I�'�.��1#4���n`a���u�j�Lv��"�!9���)��K7��~�ͬ���aU�f�*x�ݘ�w�
Wb��QV�G�)a	�Y������3��+|"܆~���Ol�3W� �$j���ă]p�Mi}���ﴟ��ޔ6.U�U2
���q�X]�(&��3�<�kp+�]��=@�[�x�"�u&�"g����/�-Փw!���_' z��4N����kh1��M���PK���7�8��^�=�}u-���/-����y���o�t:���1ιlVf���;�,��;�"�o�0�=�C�o.��D9}�T_L�L��gߏ��^��:Sz�}ɼDR���N����S<`P�ٗ3J�W��N!�!oc�������^�"��"��G�������",�	x�cK�
��_�Iȶ�6?�?�C�W�C�K��#�Cr�U�9���k��+)=��އ+�a+�^K�Mg��f�Y�6>/)v��@�"^E���������"�)_��J��\��'��g�,@�[F�f�P1nz��}+��d�м�}&B���
��l�X���	>��п����#�����
e"�� 7���7SQL��_�l7�&�:^� �ǻ�Eٔ���# Ɗ���Ef!�!���׻xdu��)���딿����+�Vؓ�$�Zi�&`�z^�ش��
��U��(+�교N��]z	&�&抢+�R�2j��^�ӧ�ԌWH=X�zcS,T�pl:�m��s��%B�͇ʮ�f�.��Fl6c��L�GMR.�;��"���s�ǣ��5!FX��қ��i��j3�\����d34�����R����+��Tbw4Es�:[p��U��I7���C�F]�����R�� ������2"�F ����5�tSq&-��,����[kn��d�E�u�7��׼�7���G����
�W����w��|�BfN`!���X�#=��v�iw`���k J�^fS��e�ܽ�Z�q��F&�����ґ�
N�q���~s���y���2s�Z��L8&>�?�ż��~�a�P'���z�6�� E��il/�sȒ�Vw��;be? ڤ��?������$��u�F.�0�^Y�#�]�1'"��*]�rM��~x@��Մ�����G._s���МU�sJ���`p(n���ܥ=���x�S$����D)�I�^~�zbqa5gR>҂>YI�/�s�:%�Y�����gﲉ��1�]��.#hX+���l�ݢ��4��&Äf%���@�5Q}FӍ M�D�D�&�L�U�d�J�����P�����X��a9��O�zI���qTi�p)�{�$G�s�0������?�K)���L�
�\�m<#��˂�b�W�PG���rW&�[�
@�~,ؙ�!?�/dX���_�^�@T�?z�Au=�o�E��ag[�>�<���׵=.w�S
�ZgU.���D%�$`�7�1 �;'��\�y���L�X<�&��b� o6��O{�r��������;<O>�%�����GÔ���& Ь���?3�&<�uevr��x����`v�_��l�S�*�����^�82�:�_���2E��O�ם�N�,7"OD;��툿�}
��ޕ6~����R׈Li��Ai}~�O�i���3C���p���ދK69o��m7�|k�%�_0�¤¢[��x2�r��g�x�d,0K˧�h�H#pI���Ǣ%������0p��<y;Ȭ�z�y̬b>�;��$�u%�6���.��Wŧ��o���	�k�q�$5_]��H���ׯsͺ��Mn%�5���b�<�ި
��K���m��ئ�������1L�y*� Ѿ����zS������Y��q&�B���}�`��p.e �0N�oW5\�v<��K(}=�Q �|��o�p�.�
w;�Һ}Qs�%�z����w�͚��x�!!��r{R��K����1?���t���?��o���R��?�s��B�9;�9�l�`OQ����LA��,	&{�_�2�a�G��i o�C=qؚ�C�|Ձ1�w)������?���^cKY�����Y�\I�tT]���GI@B������W���'�,B�[9I�q�V��0A�&LS�!�U8�&�+B:U��o��������]��Mݽ���`��q�ĥoԺUi�}�۞�v��= Ӓ	Z�hՑ� s�H� xPARq��9��
������9w�v��)2b���-5������(%�XY�w�PV V���[]U�Ꮂ��_�u��?�ib6@n;\��m�㧬�Tv�}�d��}����]���4�̦a���\*�TT"@ua��R�`3eA��H�-�OY�R�o�H��Aa��G��^mW��qy.�s��������hiWܫ]��7ؠ�)��q���Ǎ�6�B�B�k�Z�ϱY��,(�����p�/[��d��x��~v�
�u�2�k.��z��:���ʖ(N���+;�d�-�G�8r+�<��D���ւ�$N���`ȎHE�p��z�l���e���vZ�94����ؠ"��]_"R��|��ǂ�����o$M77+|%Z���Q2x}ډ+-��f��	j����z@P�
�氐+P}�&���N�©qFrZ;��̀��0l�6����Y�r@a�[M�!�����O�S������������i�Ò�&1R���%W*e��i�^V,���
��%�%w�_�)�% �؂4�0�GCs�i4i}�ۇ=0U%=V�ƈ�L�>�܌�2�2�m6vې��
M[]�3�ܗ��M�ےI��o9��I��Bbzmn����=O�7d�w�[i���^��7>�ò����`���+δ?:��a�#Oǐ���M�jcq�Y�������9彵)����3ׇT��s�+�O����ڬ%��<�>8(+�O�'��o��&��2#Ï^��L|� ��p%���4HM�"��9eh(����Iɍ���6���2�5��2�zzϱ���E��Q2��=25���5�����g,�G���R����rj���Y�A�ju�ؓ�tQ��i��mV��E�Z��z�"��?b���~3���������vu�aN��y�Wڹf��WQK�ӷ�j�n�X��h��dz�� �v�p8��dmUZC���=����Vo� ���w*&1���d�+�;i��r��7^��h���S���]SZR7&Xo~�6a/."��e:L˘�6�q�$l���I/�K"9��CgR�&,q���Κ坥�:����7�.U� >d��BWi���j�����6�(��C$�վbg��=���>�	��vg�R�W��R���Cc��JOC��ѷ�g�5�5�H���o�e��Xi�R:����<l��߈��HMN��h�U c�$.]���g�JҦG�O�����24s��q�u�&F5P��'����Y7t� �ӄ��Ig�	�j����-O�ٗ0��U��{�Q�B�Z&8ȿ���>���@�u�Ҵ�n���!=3�����dc�����D�����]�=��Hu���MT8~Fe�/g�f	=��o�E�`,! )�m�o94-�v �@�h��M	O<[���x��� ���M�9�X'��ʍ�r��/:�(kLe���5(�ˎ�|��c�|�{ ��ɸh��4�&&^-[��}���IC��މ݊�3��.����_�����7fZ.2��~�����[����i�=���������3�&#��3��n�)KX���lcD�9g��>���#�!T�ؗ;�2`�4��?�=�������9</��� ��o8�\Ο�H3M�A;u"z�D� 
��0FmE,Q��[ɻm�f�0Jvd@$/]&!�+���/��.ՙg�z�cһ�Z�/�r k}=1�C*��ѡ�T���l
�b�V���i�*��jH}ߏc6�Wcd����b�#�#S�ֺ$���%K}����bŘUl]�U�t��N�ZF��N��~|_1�P�mt����>�4g�Л��54-Mny�~��e�( '_<O-Xd9_x.9]゗�N5
�e�x�ç��Q��?�鱰�o��� qM�N"��I9��1�΂~GQ�6^��*����.��CU4"��E�H���݃�����O��c�ZKPkk�D�Q��������G|K�pX���,	*�܇L���v=dA�ID��.����k��>]�̛��1�L��W1� �mT!s�����$�v�(��\�@�ʽ+|�t��
����( ^T���w$�����.����w��tj�L�ӂ_�� ݳ8v�Y�����q��ę�y1>�E�Q8�B��������+����@:�Sg�he���k?C���ʞ :Z�/(�߭�͸H`��5���Y���n������>��D�k��>�t�E��y<�S�n�~��[��N����,�aD�h�Y�Dݐ��tJ�bBq�!8�%z�
]�h���v��g��k�S�ิ{=�6:/��Z�>`�1u[�� �ā$��1Иzj2�^7���nW2/������H��DHW5��m���4�N(�>2���mT����q��t �uBvThD�̌�LF�l?en4�*;!��������u*��|�Tݨ[j�YYaA	��#��XCWb�y�y�f;��K�U@�Z�
���Z�Гs�����QsIE�K�ͼ,d e�,��bqO��Ҽ� �c�+����UK�5^%N�v�l�*6����Qm�n�����@0�k>hh���%�]�x�򰑩���U�k ���?$����Lwq-
�\kg�����3�˺�P�<�b��xt���+%�Z\u�>4Ϲ8��~5ע���ġx��b𓴖�v^�$d�=��1��J��bq.�7;�X���^��Z{�0kS��n��R��&%%4�-|�ҍO�9�,�M�����1!�;���lt�MLo�a�s	�����%Á�nl���������s��}Y+�꒖������׵��J�0��ӿdv}�E4�@�&�,�"�[:÷sN_��v�8�ɥ���٪@���1�A���<����p\B��w��k����x���������JW� �~�{.���X\(��*���YҪ�v�'=v��}{���1+�>��$��d�0��.�s���Wˢ�>�Ҹ�X����^*w^X�-Գ�s�+m�&�����s���Z�Tb\�MFX]<�2�*��wUt�$�!����s�s7Ok����������*<��v¼�d�wa�6J`���\�v�4W&�R#=8.#�+N�a��		Z�v�y(�{��;ϝY(v#�	���3+�
lZ��q�aiW��F�3��Z���CH�g�"C*[Z�Rks�i�iVw]�>��j����l%�&��^Q�p���wo��p�~o?��{[��O����s�o;�<�4�B�L�P�(�D%B8I((<-I�D�ݸs �m3I�N$��HөD�7�^KV"�
WY��
g����O#�Tx�Y�0�\U�����{II�6;(V��H����p�&���r^<�����G.Vwr��$p3�w��E�f�i�*�_8�:ͬ�{զ����jD>���<�8�I�Nq+�+CvȘ�vC��<��'��-�t���ď��Z06=�YNA�0) {��T�l7������Vo�g�=-�0�s0}"����op=�an"���Õ���{p�/B|�Z��{	V[��N�</O��+�U���Zd ��K���Z�`��^J"��?O��T¦��xQtؒ� ��(���Uy�:�V�����jlȭ��VOd�)t�G��c������xK�����3�c�ל��"Gё�s:6��7�p��fB��2���Se�v�MC�y+�49��Z>H��S)8���װ\��&Q,��õ���¶4�Y�lε"�t<2'1J5*M����q����!1X|��)���
S�-�*x��5R��$*%���+{<�~���q����}L��_��,w������
X�g�9��>�5]⺴��כ�4��]�U}�)�����@0o2ɸ����t\���w�f�גE��@i��6��_#l�[��A�H`�]�7�y|�5}r7��-!�K������!J��##�],�g�:����N"6��]���s������J��ع���J�oD��#:s:B�&�,������� ��X4$�ܾVj,Ӧm�^�ukP����n���,�Z)�	��%7�ԓz�V��?٭�@�ޭ�s�C�ŃI˝��;Ϥj3l���̆�j?� ݮ�nD��L=�g�u$�F�$��d�͸,���+�Z��Y��6<��~��Oĝ�O�\W#�� k"9��v�y9J���E��CH\*�R<����81�c�7�ǌ)�d�^�wX�B���ͩPT[c2�$��'T��ɚ�j\�����QFc08fb��N�l��%�!n�����^�-�7��mvz�ʰ��Mq`~���fhk� h�&y{��R�Pat��5���9� �z�:��ܣ�L�4$X�#!-����������"�h�y�t����P�p6?d���Ǟtt� +J_�hj��e���'��ޥ:'ߤxء����2#�a���=��	k|k�)dZJ����aA��;۾�M ��ۄ��/拞��B�e��,��7�GoW)��HP|9"Ө��s���[+/����0���ݚ5o\�� �Kw�W��9�W ,�b�q'�"�m�)�up
�g�����ej.6�ϼA%�W8� ���$p�:4e��(>�� F�2�P �����	z�e����U�����R׈ꠇ�3�g�{>�6L�&�B7F����!����@OP�_<g�k ��9Mݽ\��w�E>}����^_#F�=�T9i�!���Q�<�����4��ߕ�x�f�2xz�;���f�z9�ݦ&g��a�Bۣy;	Ǘ9���k�؛/�I
�4��Ѿ�Y,�Ŧ�	AW��k��{�΍�E��uBuQ�Z3$���&'*LS�� ��B=�qh����2/6�#'�}�4�p��7'i�I��a]��d���U՛W�<^�vS���-�6���O�w*.)* d����gL;�#|u-�EN3���Iς����;�T� �ɺ�7��������D���i�Hf1O�+�z"D�+m��e�����'H���I��%V�x[����.X�������ӱ��o1��Wa8M�6a1nϓ��Go��F|����;�� �#J.��M>8�ա��W�"�!���i�H�����f�N�0����$����H������j��'��Qk�/�0����1��^w�r���{:ļ��@p�gI`z��^�R�\�DڕUy�s�]><���z5Car�JAI� �\��g����F]?�
#$)�Oi�fy�L_j���xtYU#-T�?՟@x�ŕ�ZO��Ul��YOV�d_��ߗ�6�N�]i�}��h�fa����5���E�v�E�I[;IȁgG��j�:�����Yy�})�`J�Ca�D�_�֝n�&��G)��D��a��@�<z�]xXlxVHYEB    fa00    1340�6Ad�C����Jj/�+1!��t�<�?���=�� �v�r��i#�z���܇�$�x���`ka�X4�/!VR% ]��"8n0��1x��ډ�A�����)Zq�Zl���-$�j"�&Q��t���7"#G-��7����,����4n��P?'[��Lti��\�]��z�����hl�+�^�]Fu�1GxUi�@���5�ᾰ����a)�>}U��f�Y1z�B��@S� ����AB%>��V)�V���vT�Km"��nЊp2QK�4�=_P��)_֔��Ej��H�>b��d������_���hpn%U�<���9�fr�cF|��:Ew��]` K��¹E��l��D�&��Ⱦ� K��|x�^�C�|O<&
N�]Ki�7�{��cj��H1q��ar��Q�Fx�H��)]�̽S.��>w)0f�s�X�wM���-cʱ;��r����{�o�k�&Y�����X�5J�q�GO�T�*}�V"�d\ը���H$$��/�\�Ro4[�[ Ff^|;V=Oj��:�׍�GVm��3MW��WU7�%����a6Nv�A����NhyJ���4ʔɟ����{��rj�Ċ6b�ĂB����k��R�Bc*�Or��I�p~�f�G�I ���O-�4h��^��Y�ֶRP��?��n�"���
�Dԓ�Kac�c�l�.o!5lp��V�
��^���&���zKֵ�)ZI�F����M��c({k�!]b[����0��<Z��N�+]F���p��{A��6��.�e���HLț��W��jdky`�30J9侬n�����?����ze��Y�
�l��L�ٲt��k����ʓck:̈,̌�٨��'֭Z��W�3�d�|�ɘj����d4���}p7�@������:h�v-��2sN�W�q���2xr��ji#�:S4��e��0K��k@4� ��k�/�Kܞ�5E��2o~S3��#LX�gY�]�c\�i�����*����F��ϕs��ɏ�Y� x�����7[a�nG������'��5�����Z�3ɒ�Y���w��*�kđ��(?�,Oq;�6'i�P{̊�����川��<o&�Q�N���G����{f��&���f.�%�_��>)�'�Cuח�
;c��_ވ�����%�y|�V���$h@plq��O�ѧ-u�G�"1��I��=ay	+	���B��&v�)�\�+{�4u�7�G,��na��B&�O�E��9Z��
yZ�������ϛ������	8zĈ�a��hݷrTqG��0�-��V�=�r�+_�F:�#�������:�9 �,�^v�'�#���2��MxzF�ᇙ{hK#Z�4 	d>M7З�B�j��n��I�g�κ�_7�0�}�����PuiC"�d�Q1���ۻ�����S�[q<=��ʽVs������x�x�a|�)�02�h�z�U��D���[w������5O��I�뼠��eG��k�L7}hM"�D�٬$�>79|��Ru�Ų���<��*#��S�u-�Ive��< �����Ek�aya����_i)��X:YB�1t�:P�ȍ8hX�Yѿ���c�5��c�	�t�5D`�7A���iy���;�\���S9κ�LҢeW1�	��ˁ�Y#��*�$��3�:����X�ޡ{h鰨���!"�y@<�5�ߖ��x$��6[?�Z2(�=()ON���! ;�GJ�|BKt�m-��r���ᠼ:�Ĺ6��]M����k��۱��d�w�##�\,a�����ԢN�=/��f.�y���,�~���3���p��&���N��	�:81=%��y��X8��j��jp��z���m�{�'��crC9{f<�C�rI.��K�j	��@��<����U�0|�1H\.�{��"敷W8�#��-+C=��	{6َEG�eXh�ɐ��u+��+�^��{Z<��a�+���a��FZL���-�b	��;�ׁ ��1s��������Ӂ�\mO�$^� ��o�q���B�����P80�/��KL~��.�qm�&3�1:�)�4��x'�T�#�(_Zx���#
�z�8���e��`�s�[E4�u�Z1������Q}� �D�������~s�@A����t���-D�4=���m7c�[���s��6�&�x�)�`	Ϩ��k�CV�����]&�G��������h7��$V�`�b���h�!P��b6YEU�nO�p�5:^Hƌ��:�֘�y�}T`��
���^?�e�up��+x�P�[A ����T������oin����ث��5��^;������>p�O�����_�<�H ��jC�"E�LHO��zz���\���f�A�e&?���4��grS?aF^\#e�7�UȈ�`HG�Ѥ^�t"��g��q��um�X4G>�ｓB��0�ư֠�tq��̻�>H����aث�< G@el-��F����@'eK�(~s�MH�Z���D�je� M7�>Ƨ���M�r�V����5'ZW��<���2rŧQ9�;Y�$�ff݉�-IpV8Ve>���厤��y?,aJ�,ks�y~W0V�k(�wge�pG�(�Sq9Mp/^^��>:P�ߘ�oJ��߬$�)����/QQy��`�׫�_��^����ݚ������c���ڴ�^�c�CYմ��O6$g�Nȡ��k��D���e
�B�h-E%w�^f8ŷP(
��V�����X�޽�J�Z�����v��|��Y�s�2���-�Nt��f�Z�|v�<�2�(�]����m�<.��^yfۛ}�@�yA�T�����^��Ge��-�B�=m_���RY} �%M��J-mfC���W�͏ЦQ0���.�.6���M�7n!�m�W����K�.2k���<��鈆�rOV�o��X��i�?�]���A�eʼ�� ȩ�'w��	�Sa8"���1��d#w�)��+�6���ho��0��(3��庰���Y���+>��U�PC ʌm��R�wE'g���I_-zk�O�h����)߁����7kQI�W{�� 0x����u(�Q�~�}�꾧�a��L���X��(E�{�],�0�O �Ϛ뛈��[��Wx�A�:Ŗ�D�t������P+�<2�&P�?��) 
���*u�my��H��ۍs�@��0�T�L�9�*�d�j�`�ymg鼒�MӤ?�vl}
��(��Z?�R:h�U�5W/��h� ��[oϊ�5�)��^�*�D߯l|
1�l�3.b��H�O �S��L1�:nY��F{K�+1��3���x~@�=t%��wX��.%�y\y���jZ�/�-f�SPb�������ԅ4;��I�A�Q���h��&�¢�Xm��-� ��'�%g9D����9㫺%>�O]?������< ܈?�t�לfxbp�В#���[V������Z����[����4Mh�+�i�0��hc3/����*����N��#O0cJ_�J����]te&eU���f%wQ]K�6�⵷Î���*�#� �gםc�'�|�mV 4cQrx�:XH?$�Y�c�j�K��!'���� ��&%M�{N.P�^3g.I����Tl� ���П��%X��p��@�bq,N�x+?Q��j���%���9�n�5�)�L�x�EoQb�J��*cw�z[���5�o�cZ{(8�i��ޝ���yJA���c��3¸R�����a��զ�PN͖ނvk*(��rp�\����0��ho�kͅK ��1a��w]"cVc�Ɋ�~z��.I����5��X?i�g Έ�����gM�P�����UȊ'3�iVFB}�^�7"7��f}�!m����H�D��{�؈�J(�:E��J!�x�������O��.J~&Q=&?ă���H'������U��6�N>@V�deF�/��6bj��w4[��c/uP�O���R1�}�m���
|�~n��_l �35��Y� Q�*&�T���ߘ������4����n�7�Y֋���3'w�g�i�,�>��������Y�^ڈ�v���8!�ư���ᏥC>^n��	ۿ�S�7�l� �|�K��ne�WШ�@W�ho֖�*~���6����������(�[��IЌ�@�h��qʐ73D��s���~b�d���]�h�皮�Őb���a�����ޛ�G�S*0PĠ��ݫ#�c
N"Om�ꯝK�^Ĕ��bצɗ91Fh[�/7ˍ(���p��E�f�U������n(��
���B}^FX/�:Oeo�h�!�
vM%؟K���y��/�0���+'���S���5�I�����@���9����A�� �c�Fر���MEd�˻���P�1՗�ʰ_Y���2>�EӶ˂�v��|��`k��J�-��7�AxM&S_���2�j=��N��&/�v	�g��%�.��?K�Z���_���/�T��^�_ӡ�M��Iu<�*%��HR�P���ͥ��E�Ht�j�"�w���u�]2L2�uq!3�K$�#�33(ì_U��Q����<��uW� ����z z��}"���5~�!����r>a�>��>�O�ڶ\0Z��W�b��o�@"��嵪c�,�!-O\�(�̣s����{��;Ǧ��^a��n��p�݇	�1��1/BB4wb'�B ~������'+��t���!<A;#���e�F������V�uU+���x�|z,'2\�2߁o\ށ���5A�a�X�e��s�cF�CMOlJ��Ky8U}��m���-2qE UxȾ.H��i��x�&�I���a��ք�t	��YK/}�Z�n6;���%XlxVHYEB      fc      b0��l;��K_�te�2�3�x�������>�U�J�4[���,�g'-�`>8M6 �l�}��+�� �"�̖�I���K�N
����3U�g
��R&'d=��2�	�I85͹�ߪ;��H~*��O���h�!k�gn�S�؊?d�Ӎ+�ę��[]��z��;�̜L