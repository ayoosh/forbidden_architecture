XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6O[ؿ1���'A�s�=�j����vʧ,ـ�����L��ס5��"�d��]6X��'�x���=M�v��@)/)�h� �z��5�j]�!!���kLWD��	�P����d��t�U�Hlf~	P�8[ӀT{��om�8:��徣���,ґԁ��Sq�M��o��z�(w���/^}?N:������`�-���z����M�g�L�~�'�o�w<�0Pu>?ξ���.e'��˴�`n��i����tx�0��*N�X�YY��1�I��c�K��MWt�\E�]����"���/�@[��"��<�W@N��IY]�G�
.����^�����
2m��H"��م�`y��(��R���L�d���7�F�X���"���Ϳc��ҀS@|��-����#	���������G����c�9L'��7n�02�áfE������A��<��{!v�W����|�ǯ�$�2�4���>7�ڐo���%����Y��F�!����Uv`�����y�!+�~Ŕ������n�%��cG쉰0���52�F�����w�.\�B�rsbG������
<�i�:ulc.u��Q⮵n��`x��ik�.&_��#���*@�_� ,AD��o�o4�&z��7�Q������Y���H��Ƕ�ea���x���~)�*���������������F+�nD���	h�	�N�<vG�@�$��&�k���j ����>�7a��0�iC���w�g��B����<�J��7�	j�XlxVHYEB    aa52    13d0�[����kQg!޽�'#�7����&��k��J4�ok�j6�bp2�.�#)9qP�c��eJIR���?��CA�%����E��d��i^�L�Z�d[���P�#F� 4h��I��_��hLe����z���I��A_���x����z.�9���"C-ʠB��y�Z��P�h}ؠnÙ;���#J���n���t`R������ŧ82��8]ׄ�g��tw��߁��6��	���a�͍ᱯ�P���r�{�fLh*4ynkӤ�s^��q�%��MQ����M�e��8��]j}�+�\����<�zAf7ʫgɧ_�$x�� ?�1p��Y7�������W5�(���j�p� ����4�<�#J� �qe��B2e�ro�����=h���;��Yw
�-�h�����,���ND��:��%�VdlזJ�	R��a�h��D5��[.�&��ۣ2�
��Ԧf�;8���v�I��i�+"B˽�\[�ͦ%���-�Bط�Ց��N�V�[�p_�;�1b6���CX"b#X~�ͅ��ì��x�W_��ʈ���HȀ5�ҷ͛��j.�����k{��sF�C��j2>G�R���i*^E�n�{Ş,������n"�u�#�K��KNu�H!���K�&r:ud@���`�����w��jH\:#I%]ǒ�:�w�M�����U5uloÆ׌�n:�YXԝ5�(z!��w�'Yۗ�G�_7'X�r��d�3�y��X=��WZV�܌D���m�ޕ����Y/P��V���[:LQ�@�!�y�4mw̌��cz�fR���4:F8s�u��N@�.����(��!w�&㠙�3��:�NBڭ:i��[\��!�|f}���*�������?;��	�'W�&�㤎�[���p1��Bq��m��/��|��1��ړ'��A5�D�������:Z����ft�B�P�t1�݌Iқ��nz}��P7��@#6���q$�#�2�:��-0�ֽܥ'��HqJ�Z�#��J.�;�'�N?i���	���n�a�s��\��Շ�]�a<;x:��g�L����|n��_c¯!�ya��RG�_���p�ES��k�ݩQZ���P�b�5��x�����z��|8퐿��B�x��Tj� ��&�� 85�t{�>k�)_J�<��+civ6E���� �M�P�! W(,�޿��wY��MIy �{�>�fn�E�|a��A˗�a�3~:-�y]�'��Q_�#�m5���1VQ>U�a�և��
:�1�n����:.�� ����� �70I�ٷ�|w�*�ЦW�06[��0���f|n����7?Ug�9�T`��St��p;�us�z]s)�\�O
v�9��[��Y�5���&��d���8$�?�B�9)A�Q�&;a�!!��GFUzHU��h�_��XB=�qe��`�0�K�W�F
�iJJ���}g�gk$9��(�����C�Zw�d��%�^: �tr%���S2�H�y_mVդ��Ʊ��P�K|� k"J�:�� M�BA�q�rk
�����B�T�uں�%���!;زa� �8�e�J��9w�>:���N醤n���d>���[0���SnU�/��]i�Ū��c�b�4�V��G|�s�<ÆH���&L�@�H/Kt�7�쌤�+ecw��"����
���ANH��֏�h9��^�|�^�RR"Ny�.�h!A�(����z�4�7P����p",LT�5��"���^䫳�9S����Q�l�:@�'m�� W�ý&��⠹_���nW�n �k����#G�l�)��HȶN�y%���p`[�F�~�<�y�V�����,���#s�U8�M����nM����>F���A�dT�[��!�?-
K�5>&u��zz��:�N�k!�(ш�_�r[�����{�ϠDu��u�������E���*��5�1OP!Rh> ��r5Xp�1�n6����tH�6���u(� wD9���H#�/,�����#C&�}�x�p3��8����l���f5v@W'
-%��'0���U_�~v��"�S��φX%|/���i#;�@���X:�?�Ρ��_�UY��	Ug����c�-<���;I��,.|�@��T�����È�A������s��G�ZpZ4h��L'+G�x�)�^��O�n֪Ŧ�V��m��5�|���(�D�^����/��D�jX4��X�7 ����2?��"�3i�(�"�E������I�/���AF�R%s���W�.w��c�������s$������t��f[��CԪ��|�E	�?b߭�5p�h
��J@�V��}M�~5\d�C�� ��_*xt��n�U��
�	�2���$�g�uv#��K�����SС��!�1�>�}�0�c#dv^�u�:H��6����ˇ��1ܽ��y�������:F�dM<���yVC������s=I�v�V�;Ω�II�Y?�������9T��W&�ڪ��T�D�v�u��i��$2�89�&[0B���	2Jd��d����Ş�?�Lp����7�OX���|o9�rԡy׶�ap�C���08l�`:�)�9j,M#V����EL��ţM��;i�ɬ�#�ϸ�'1�aQ(��آ�V�o�׉�uk����f��ѷ�B� �VӺL���*VT�4o+���N@Ye�i5��1�H��ǻ����a���O�z7K[�k�=t�KV�6�!��n����,���o�'�|�C�\�V�f�S��z�����d
80�!�� ��=֟Y'���̡ge��"���ܻ�������lm��r�W,^���F��.U�
�V-,�#m�P�|N=lõ���C����?�5qBb���F�rY�t?�_a��n�V��2l`��@u:��/4j���P� ����lh=��q�����[rV��9��3��=�'+��Ǯ��=����'k��?���9qrp�VT/*�) /(ޫ�h?���-ˏ�p�[,�8ħ�F������Q�h�MK����0��� ܢk!����C�{�2#�^�H�/I3ȲK�[�x̸��q�pB��.��r��u+�����o�1'~q��[,�����"�.F����=��G7!�|XiC�3T�Й���_�9C�R��t{H'��v�;}��	]1��p}��w��yN�Iu���iT�F�X21O�ʵi�v��2�
Jd+�����'V�с��r�G��EI���D���� q�	������o��Mdj/�~/J{�<��X�Q�;��ۏ^+�Z��-dG�Gx�,˳���g�����1,?:W,�<ٚL�A*�����R@fX+�����_%Kv����NT����J�:m�}�Y9G�E��5�+���aKy�"�*讞���K&��ޖ���g��Rع����L�x�M _�i�x�J',Y�ُZd�Ӻ7��V�����l�0Vr��/���W�Bt-�߭õ_i�C�I�.
�n��N\Ðf# '��_���n���eO~��ic7!S�4��RS��p3H! <�7�Zqo�{���Vl*���n����2S� ��ɳ��`�&)V�,l�Z@�N�Ѽ���SG��~��}Ԥ��� 㛥D�RC���ZR:����̔um���↤,��L�8�0�<�2���ܭNQ܀­��wHN��@�׎C�׿x q��M.�`?d]e�R��՘��Q�iZ�4���v��v��q��,�)x����!��u�
IH!M!2��rF2���|��R׍�K�.b��A�h7� ��T�&tU�r_�&���»��k�;�:�<?Wr8��+�f�r�F��Le�7��1�%���R�"��b����C��k�d�m���h�w��>	w��E���H�W�h���,}����m~r�7oS+R珼O;I4��ԟ�D�����X�@�S"o+s�xC�趑��
=M0��	���C��?��+��Ȯ���b#,�]�+^6a��)�";UDطTdoCrN7�fL>���L��QQ�c^]�UaK��l;�m����~)�mKkh��f�(���'\����\{�_��o�5cc�8I�]��+��[Fh��� ̀�E�b|�����;۴�`�p�:`ޢ�B|�ID@��:�4,8��#M2���MP7i�vD^��؛��Ҵ��h.eJ(EC�<Xu*$#�� �m2P��<U��g���m�������,C�1|��� �D�)���f�c�XL7rژ��X�l��%�Ï�.P4G�,�.�Z56Z����G�jM�=�ÿ�v7���Ө�F� �&&�d�W��;:�pL8��P�zK�]���Ҫ=�f�-R�����b������）Q���9�	�Q؏G��nF$���M�g�!�:����Iu�HN�AE+����A��5E�|o�%��`��vY(I�W��e�2'�����\�|7���:*U_&I��ҵ�H����C:l��B�BCCYcY�h�^F;�(��3V��7p�Ct����g�P�L���NBD/(f�C���:��V�-բ�-�]��if�RE���Jlz�v1O�F�᜙���N��z�1Ld�	9/uA��UN:\ݸ���#k�<1x�ڭ��]��] <N��ߚ!fF���#<M����I����q���*��N�+_��{rV�u��3��r�J�v���B�&P�6�eO�L����Y��8�(���t�װ��tKƃ=,�DH�^TK�Ў��
��a�w&��;��L$7�b���]P:��z$�~;�S�Y���<�/����`X����$D(�qn�q�گ��e��5F�e�N��KyAw�R���P#�	��Y�]?�X;����jV���/$3��˯�Mp�����9Rs�m[`p��W�Y���؛�70�h���f-�bO���	-�%����y�0�b��z�!xY7��ښ�I���+37zj�����S-���x���|E����&��4�?