XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z�:c@�dHf�
'�ܮ������\�p�s<]vi6�|/��*��ٯ+}�o��d�8����_Q�/y�y�Ñ,qp",�l��y�4�J��w�"tT(����(�iN�`��MU����Z��Ml�ܫ]|�|��M�M�k�SBnI�#r�|��sv��G`U)��Zu]Q�Yc�j,a�a�i}) ��Zo�G�8��*�'ԛ��L2���R"���*��O�^��(�Q�l�k��s�(�pB�Tnu�d;��q���s�ta���j�0��%���y��=`�g��gd�>WMa��=u7+i�^�K���ӗJF�)��]��\*�J��U�s�R�1e�6gG��E����l?��Ƒ�D�HF}ia=J�53fN�`�&S��߹�
�����Ѵ�,%�԰��m�ܪ,w��ʐE"����	3b�TJ�f hZ*�H ����#Ok���Z>_J��qJ��6[�"v�.lhd�����γ
9~�jI�B����[We�D�����L�e]YlL������Ӑ��S�t�#���uz���y�ʎ��@v\�䑞r��rT�Zz-��&�t�솀35	k��P�9�n1wq}�z�\�ț�QF�o�)����9��^B��`ǝRU�x� ��zÎLK�=ly�������ψ>J*Y�`)V}���N($p���早�wr�C��ޤƾ���E�!����v _���;QJ�f�y�B�j�&�~i�^_eq�8i|�9)c��m�{�dDZ���W:XlxVHYEB    29da     af0�b!�������f����W��@�|L	�!�	X>�Ku_ُ�MS10R� �H�Q×۲-�����웯-:9D:��N���$e�aW��GCM�#����s�9�� :ǧ��+Z�gw�}���{-�D�<��K���C$�_�Y�th�"����j�f���o�/�߉Nr\׌�*�A���?` ����D�T��Yop���N�0�XD	o���"�$E!i\Z�xF.R������-a4�0.�_��O��>L���e����ɟ���d� ,y��p,���悝�Y���U-H93������k��49�&��'J/ #%U���aɼ���l�y�	"�gtQ�&��7���SڹK°mQ�pzP����+`{D� -�H&�E�p��{�|�e�=�ȵ��a؞�`��?�4�9<Y1Z+�������>M#���ޅ����f�Z^Ww^܍E�M�K�r,>���l3][:��'�w
�B"^. ����B������ �1��T�Y1^�j%�KY<�d�	ށ�A�(�F?�/q�)�%ȕV(�m|}')y�b��<����xqx�ԥ�f�509��^�Wm�J��6�|�*>�����0�L�.��j��-�zliJO���$��i�EZK��M�����R����s�t� 8.�V��/�ʴ6ڥ�!��� ���w�{�id�P#ȣ�u���v���aˋ��?�`t�Ykn֍bN�b��<����d1^	��I���� ��1���c����:+遉,�#M�	o��w�M�+&���`v�Oo��\�)��ƳX��?�"��e��5�=�)Ԫ���z��E�&�XpJ��?�Gϵ�E3���.�܌�5�:��l�L��a͟>c/�`��~� �'���J�r�ܚ�f$�IW�I�'n+�ή�?|G108�����o��)0o�sJ���B��nn�ܛ��]'�����'���N�y�M�&�:������W;���:���ϳ��zV�/�h3��Ii&��0%����Q�SIЩ��C�^�TR=��j���G}��	��IK�_>�՜�(�¹ۙ-LL V�X��n'���Б�)��y����t�E�AՀ�
��1����ʰJVr��=�Ѻ���nɠ���'�^~( 5�I�o�R$6hg0���,�5��A1�7L�( e�5��1�ksY��[�mZ�n���^Kޮ@CR���9�u玟=2�eo�"��l���>��N��|�ʶCİ��>1\���B�+0#q?�:q�\��eQ1��K�z��!gtś2W�Ɗ��l���ʙ�=m̥�h�M�.I�'�R���c�r����l�3�	U o���ݞl�(�o7N�t_��ro?s��e]��qc��(ܳ�=G�I DPa���m"�:%Ϭ��wn���s5��8����Rw���~͎��k"]p�|mJ:S�-��^�p����� ���p�4�UV��-w�E)2����:�����Z�iX�Te(�F���	�	K�"O�9_�?��OQ35Y�#N���#A�Y��3$G�T)��4e�pG��co|�l�YF�|��.�֮�ے�� T���3��>��H�~�ʐ|֗�|դ�],q�9g9��l灌�j�%��P���""��Q0��Ζ�X_KV�]/V��Qs�	s7D���I�\����ܓ�Y��X)��G23�;�ZX�E&X/�|z�qg�P)�)��B#���*�rc��oVi���hDygL��X)��%c� ,�m�i���p�B��Ǟk(�<eMPKIP�����0g=��[�>��^���ǭB�˩R��W�oj�b�Ām�U��yB>�I�*��+QG5s:�4k���~|�6���	/�'�n@�-X��a�΁�j����s)�J��ُp�{\���
�MP��Ĩ�?5��,
@!L0#&RS��[g99!�zO�[�/Չ�b�0�.]70IJϘf�A�-��omX��b%,���"Sd`��v���T�9f���߁Ӫ�Y����F�D�af�^)�r���$��	ֹx���p��ɤ M>f�i��Ҥ�H�N֛���G��d�W?�.�I��v½��t� ��x�;���
h�ƹ�iB��VUnr�|��zI�K��C}���\��l��LM���ty�xp��#'�q|��xa1�8hX���&�Bd�eđ�~��b�uJ�G�1����1޳���bB�׷�^����ϒy�Z������Y4�X��B&�Υ���v��Gs��r{"��C�(쫛{x'e�cz;��o��7�g"��<xÛ��	
Yָ��l,�{ҿ�g0���������O(����.��JH����O>�KUU�^da$�ޑ͂�<8)�b�j@q�T4��Jg������?��2�(�p�c҉��۱�N�w>b ��w��Đ`j�����Ќ:9�=n�8S��L���l�Q��H�+J��$Z����x@�1Y���kI��E�Tu�M�ϖw�>����I��<�}��!_׸���� ��!���"�+�S��s~zFN�P�(��{Y�n|��B��U�ѿK8�9u �:��!!���1���u�%
���٫�;��?��~�������gãk{F_[���o$��)�����;�;J�~!L��v�z����q�؍���g��8�*Ov��P���u=��e���@�dH!\������5�a�$�'�����t>c���$�p�_!�H��Ì��"_��x�Q?j���C�͏@7v8w�