XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���nx�vp$��q���pDD\3#�	��5a��b����Tô�^�� K�^���������N�>S�P��|,��1���T_�3�Cd���e�"����������C��'����M���S_��w'�u���n�w�|e�z�Hz�r�*��7����HW���|4U��+�P8p����� ,�CQ[=!�n�ҳt����A�(�l�S�5�W�Q��6.��<~Z�I�T�9�7w�7�n_O�g�	I/$�=�KJ��{7Y���-ӏ)-=τR�t�Pgg��|������(D�iW����"������T��8�"��%�{P�c���+�l	�������҈���V�"B ��$��h�"Xƒ�wZa��I�{�Mf6�M,������5u}Pi	a/uv>�f0�^+���� �`V�hbWڢ��#k��>��骏F���0��@�9T�4�Fj憲���ӆf���Ф�	�BH��[�}��%�$�П�w��3��(�(nfk�#e�r����a�f�%!�O����|�V�v��'�h�?D����?��X� uE������ĖDN��w��)��U�WJJ���[p��k�7
��<����.Җ�M�B�������X�5<1���L	^`�li>��r�O�D{`�T�E�������K�<(�k��v������y�yh������˞��boi���=�/;����l��-:����B�Ȥ�'�q)������j�nre��XlxVHYEB    9f13    1bf0�X�J�5���}/�W#e�X-Z��"�$!	�TB�$�l7(���=��ߞu�no:�n��!��s�0!�(a��A.gb(y�	�rCw�A��ɑ��ď��R��4��<0�?���o�5�P9��+���e<(�D�`~]���6�h���T5�p1���-�7��F�f�������R��T�2j!�����G/�(1�o=��%+Y��'u~�\r��:0����`��!�e:�E��k��ђ��m��1������w���R�q�E�DP����g�^���?�_H��͑Xh+6l�]1<�[�v�zN{'��׃�ӑ A#\vTj"�`�v��4<Z�ˁ����?�F�[4�[K�X��la���T�i浳����y�}neB�r�����.i��U��gl�ľ�ԓ�tA���ed��.���ٴ��@��H�:���-in�N�w�s)n�5eUir��o\�������QZ����"�5�Ӭ��+k!_��Tֈ0R���X��Gٸ��2q7�j�gڼ]ԓ����6Hڞo�C#�������<�C{`�g�T	6�}[�s��^j%s���F�[%���;����h�5C���vz�������ح���@U)�첡�=�'��5e�L�9���J�
����<"�mBȡ^-�Pv&;��/3�,x��Cv�DqN�P]X����-?հ�=*��3J뵣]^�خ��¡�Wv|ǐ��8Y�
.4�~",^di�������c}tu�"��+d�60_�2�_��	[�.(�j�%D!�ت(�F-�O\�Q>���_Q���("J����/���@RQ(�Y:%�Tc4����������'+,�cF�a�@Ԓ�D;GVu�+رˮ�y
m�>.�q���u�UB�_}R�n�Ͻ2w�=h��:��{"�d����asT���/�~6h7ˏ�$'��2�IˇǶ���~&?�$ڡ��w�H���x/O'���j
͑�I�/�[�t}���r��*���^$K� �]9�2EjZm=;na�-�[��+ioX�~�­��4E�!��w�W!(�|��:���>ze�\�Hs=@��a*׮t�����Үi<�\�����2xIt�Խf<D���q��؀;-@QS	��<�_�HV��`�[04��68ka��e����^l�������6o�E�ɫQB�^��^0wF�J�����
��i]�֋��/�I�#y�9�vhM�@ܬ1�Mݜz��c�8�o�(�3�l��.v���V50p�ь�P��"��zRDK%:9�+<�N���!=�Xs+
���c��ю��dƒ���4�3�i�'��\~Fn�Q���UCf�vo��H�/A��J:�0����v�!`f+C�>w��W���"
9Q́��Y�AY5$��Х���1�%}/��:��ђC%�,�� �q�z��@�� �MF/���I�Zx3����4�jE�A-�� �����!���*)�P�K>!I�[����|���}rg�h{�*R+T��׶5��Uo��%��Bֿq�]���]˰�d��I����R"w�
�*ʬU��R�&���y����w�����޿��;y����W]BA�S#q����6o��eؗ]ݵ�MN�ƫž���\	��3�U}Yz�T;ǉ�D��b�vK�rD�ѡ�i�a1��ۆU�<�%������Z}�ڪ���#χ��h|���:/(罖  �!�I��u���Ԅ?٦"xq^���By�7o�L��K����
��3���S�Y7��e���H֌qz<p�~O�\F�<i�n�^Q��`V��axB[˷��8�*���Sr'=�S�3�����p�C�DD��.�>�e��!�$xnk.�LE\`��"V�&x�D���E�S���䚬��'y���	gaVe��Ė�V��8uH�n;��MJ��@��pA}�z�8+�?]tڔ�D�e���F�҈����=�馮W3����n�,ߋ��}���!"hs��"�d� �V��-E���m�a�Z���d��k-zϲ�1Re�cǱ9z��$�6n�h��N����2�TmM�Mm[2��(�VL�:��97�s2Wg���P�B����?�X&�|�Q���/6��B�!;����4�D�S+��)r$��䅈͛�!�h�Yv������i�UU�&Yna���C��(oDD��T��B�ᩑ�y��?�B���]�������Y
��n�����l���7�t����_z�����
y:^�]�U<��B�c�r��#j��-��o��l�9�p�FYz�m�]xZ�2���D�*Ypε�ˉ$�ֈ�T�;�08���oc��[>��_^����`���2R#4[l�)��ir#����gP!�����PZ�o���4������֯�Q�Jv.�s�2#b�h�ۊ7�s^O��Oc<L�$b�`;��8�@FMo�`��8�y���
��!)F��m�Zܾ��,�0�.:��BRc1t��x�:���䋱d�,p	�֊vDN*^��2����7���3���$7��\J�t������A�_�D�x�Ԣh�<��JѾb�yL�~O�;E'�[��������1�։:�=�mW�u�I��?�=<P>�S$`�%�ً9�fx1_O���� ����uܗ����OS���; �~c�$�t(�ʒ�|N���+�@/8>U1�٘�?�],8����2Q<�#U�%P u�`�"���$�������m�mxk;��boux-�	���~؅���Tf�GbH�Q�$K@oF��9͑M-*�ֻ�[�GjQ�}w�M�KG�ֆ�,q���{�Uƌ�?�82!{�G����������,��=r����3dg�P�DF̩DZ����a�"ֳ~�b�c˧��9���_� �[��=�/'���d�8��I4��l����E��F]�Z�Q�0{��Nʴm�PI\����b
�V�5|�D!_p�q���H|Y�:�
e�Qݩ9��2��kq+K�.��?��Bzk �{x�1��M����-�ũ���Biq+��ts�0�����\@��N�T؏��夷7[t�P,��,�
�xv�9�|<��>�0���]��M��A�I,�Ǜ1�H�&3���|1����Us�r���N�|��9��7K@���@�uY����[ m��
�(C���7��\�rur�(0�1���/�����Yyng��v��;͑���b����1�MQ�]|�)1�+	�3R��Y�}���g[]�-ɑk1�>�gq=�jW�>,�[xQ��^��.,V���tY���ծ��}�ʗ�N��ضZ<�DF	�/C!}U�w�}�P­��/��͠Vj�ƪI�~Н]s����_]���n����b��x� 8Gvq�_W�!�y�C8,�6���}S���/��G�S�R#�T��+��/_u��H�@��Z9*�<����t��V�_���56�7^�`����g����Ƕû&�6G���o�tk��=R�t��axA���i�[5_��O�>���<'�Ĺk��h��s��Cc8�E�q�S�Գb<���	^���c̘�ke[+ƸtxL�(�(����3������$'�w���m)|�1Bt$�h�9��7u�]��@��0�}L��������[���\�2��c�:Ir].=�u��-��;	?hNy/r�B���H�9��hs�����\�m:}�-��x���ċ�p:��0��h&�B�� x�������LD�Tt���[��7��$�E�/��R5����IE���C��E�i"�kFou��g�і!�sN��-K�eK�	����s���O��;�?�T ���Xȋ;��n��,�p߲^f^�\RY��lI�`��X�=�︒g�pVը�Ϝ�e�p������\��S�c�\l�[��s���a���6f��#���.��z*���k��f��uŕ�[�.nf�9E��'�Nb���v�٪c8M��1�P$�J�:?�K�����M'��������{����O�(�C؍�`/�{�߄�z���
�=.�{�%��rZ՛W����4@~��s�~��Z�lƷ�x3O���]�v�Xy:����aW��Z��!��'�k�D���\4���3L�~����������Y���]r$B�3�kgZw�#B�n��!*g�;*!�<3U� Uyt(v����&��}Z_��xpg�f�^`��qs:A	�$���J"�R��ڝ�E��tA����T���'��|�����A�+ԫe��	���U���Q!�'��,!�O�;��AQo�7�>�&xCC=j��/L�B�����4��셋�3�I�J�L;�oSx�0�B	�̨��p��徴#�h#y6�x�l�MW|�{x#�9ǋhN9D �5��ހ�(`�G�M�$h����º�3��r�ß)��S��N��}��Ѷ�:S�#l�k�8�lU>��?�1�+�~��אf�Rar*�(��e�b'�l���£*"?5]z~��$�or�#��W1�s=/\d�/��>�p�OG�����RT�?���,vD���C-��;`I�:U?k�M�Kh@`�r�WS�Gk��.�v.%�#��;�x�dSU8g�65�6W���RP���Q�4��+��ݐ��'���n��ģ�X�Q�$q*"����k㊥ң��^��� ���V�dM�/���^Ƙ�P��Ƥ�`���|7� ����� �\��Mʠ���F����� lx%�g�c��I�3���kCY�PТ�(�^Z&�g�5�!�B��<��_�*7U~�}���X�<��D�,��x�D1�(E�����s���<��$��1��
K>߲Bt�cX��D��j.�n\��*���=>,kYNA)k���&����x��I"�oO��r}�gQ�&n+u};�D�n��a"Ul��r�B[ha�	��[�!�.)9׼@�8�BM O�
��p��ENl�J�yF����|=���N���l�tl,庣QI׎�6�((��+�?]��Ɋ�j���Q����|��RRײ��>K07��`Б&�l'��֓�m�6~�;Y��ƞDd��5��x�m����5����c�Պ_��m��}�m=�[aB��U�;�)�aeU��M|QB4�ɉ[� %~-72[��{ڗ�RD�է}Vޠy��M5�/��T�� ��W�wIt���	��6���i5q�Ct�A����:yH�'�1a���������{;��Н��e��Y�� +�?�+���Xx�n�*,��e55��
_S-�4��&���v����rQ�qo!h��_G�J���|�X�Α1L����BKׯ#N�N5�+��8δ��5�+��R���3
#����V���8�~��KZᯣL��%XA���7�tlU0�C���& �����F�*���/�����~��t���C-:1�SNh΁�(�W�'c�wE%�b�,Ez��s�C�;~�%N&�/�C-k��PС����L˼Ie$u;�.��u��x(����0�(����Gz���$H�[pO�����Ŕ���j��?���N����Q�H�B�� 4q�
�ط��I;H�Ū�ٞs����0�_�R��o��t�Y��s⏖��P��SQ�'�!'>U��2�$|&t��q'M
���5���Y�j�ta��s|� �c=5ciY��2>��S��cK�Ĝ@*�S)N�;7_���/)Q-��x�w}�Y�'��&B��#���YI�"�yC�b������i�K�%7�Ѷ�ҏNa���\$6���F�[s�\��������}�3..����]�#1����IrX�z�`F��O:@w쀓�
�^������ֆ��Ž~@&��4�5U�4��R��=�������a}x������$��n$���p�����ǼR��B�
y.Y\�:\��;�)��ӆx��n!H�W��ha�j+}����.���&-��OL�y��_c�'c��І#:����U�A����y08�f���D�e��v����$j�o��޷���M���f���;S���:˽�����o��|�\�O�`.�лI��O/��m�0D�RuT�@f-�ة�m����i���,��=����,����镴� S7��I;�ū�qaCn?bz��}�����OXw��z�5L�QU�Qɂ�%�9z���Wْ��e���6�z�9e��Wx�>_�慲1��J��UGti̛i��t���S���03�ࣩw���^�<Nm�,���2��bV��.�ݯ�5�}��x����@"^_��T�*�Vqnf�pG���m`�rM��(E�z��\<�h[]�U�d�Onq�����k���G�YU���2��BLc�^q���3�����5ߑ=��S���?�qɶ̒E�������D�0ℑ�l����(�"��ќ-0/�����eǚHK�Ҳ[�I4�1md����+��ԃݻ硰�yƜ�sc����˺�-<  3\H��7�X�FN0��hv4٨2��vڷ���������q׈��Iķ��k�6����6S~6W���G�u�ENd��c��㢲,��G��),�4�y��+�,���j�M�Q�ORB���rزL���
��zխ�^z@��A�T�#���N!.���s#�;B�B�O����Sp$
��\d��at+`;��9vsfn���o{�MV�����B@?����NZ���Ť��^���{��}UQ�N2��JV��i˴ y�����wr���؏.�xN����>E��}'��j��>��+B0W��^Y��jWىN�v�G����#�Q*���x�s�crx#q���Vh9��M원�դ���c~��v_�kt����8�J��X{������o������o ���Lp����5��v�E�jȯ:����P��pC���S!���D%��LN
��Z�ۣ��W�Q�ic��oyږW5F�ګ,�5�vz��mCګR
'��
�'�[�Lu��y�`�/�/���)�8��Ç������T܆����2��