XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���)]$�#��Q��(X^����Ce0}�;�� �q��h�P��_�%�"i:rR���� ��Da�R�Ү�L�E�U|]�^�ߗB.<�Lo���t��H]P�J[��p�bJG+�WHJ����in��i�Q�v�x�w���6�ދ�}�l?,���t&iD�:j2}x���L%�v�Cv��p�j&9I̽� �oIr����c5%gx+�+[��?���ލ']$~�ŕf���I�]F��6�;(�A,A�r��y�L��ȼj5Q��#���[@�oY#����0^o=�$�_.���gj��ʐ��(@�����߯���&X�B9�1BJ�k�T�Mj�������<K�BJ2d2?�
���� �����8��[�s"	�n0�ؤ��2�.�����3�=� R�]�9N�:vq�{���l35��.��i���������	���'���u��An����=I�������.!���z�7������}R@��j�k%NZ��i��9r���#�L�v�i,,?�G�(�a
v��4z�o�-�}>;�mUQgO*��$�R ������˗�F�Znf�ť�,!��֡�<N�=0��~c�sh��t���{�K��k9�J���f�dmvK�F糸@�.x`��\���EHV&�ʝɼ� �����@}���&��Ἴ3��v����p5��f���~���F��0,g�Y�V܅����	9ޫÆL�C�Lʳ�\f�e�?'ǘN�g防����ߛrH����XlxVHYEB    fa00    1ca0R���y��1;�� hV���r��|���� ����dd���u����sD=�����X+ʩ�r��
OD&��i<'���lt���#O���HO��mGY[���x35�֩Q)����� �O�a�����,�0�^�|ȱ�?�,d�;�;Wy ���D �z�8PO��$��&Q��́-�РZ;��]��i�iF�Y)(����_5��� �#��xӂ[��P�c�[�>G�=׭m�E�U�`�^���6Za>u���q$������eq��O��2�<����X�����w�N����-��\֒{�t����g�s�d�/�`��D��|�̵�X��Qٵ	��t95��j=���qt��.%ۺܼP_?������G۟�-Q�G1T�+�(u1�"|�a&\��<H;ԕ��
�ؙ���8�h�M��\�x #j���c߽���.�|굋�E��
@����;��6(F�ᥜ�}s�k��(^�������EZZ��y��(I�ϪOt��C���_�$��=6�ThZ]��ayt�+�ޗ�sJ���J�����+�B!�ʬ�`��:������ R��
}�|���^x+f�!S+���!o!�n�;$��ʠ&��TCư�ד�h�C���om*�"<����g�3���_U���\5 �C�e*��@m�Kl-��&���T���w,|v,Eٍ?x$ry0#@��E
��|�z�n��K��0�l��HN��%�JL�k
�NO<���c��LoG�C��t��}�˚}�G9LwtA�ϧP�B�B!~���Gn��o��F����[�G\)+tһ>�R �	��X����)eH<��jۜ�hV+ܒ���w�����S,C�+�=300�,��>��������>�kR��;ܼ]S��m���`���vǳ��� �\�q�C�vi��I4�Ӟ����0��֔�V_�Ck���d�^$�d���S�0EȪ��|���X�˰�b��_Q)�3������B�k#|��豔^ϥzD��c�������:�O��.���n��9P)��o�l�*=B��oɀ���:����e{u�f����O�/B�
˻�`H�'��K�'���l+���56�BZ�:����|\'@��
(��Ě�ȁ}�p����ꛔ�D���3�7:�F-Ûo�r:����|ڳE�z�@#Dq\o�y��uU f�+�0��l��#��zbb�o$�#����U��&��i\����	��H��w����a�����:���3
.1\��zud��$���n(j��Ӝ�E�3���ZvUQ��U�v�F���-`�ރM��N&{�=f�'e��C��m���M,����;��#��$� Ydqzm�1<�ܧ9=�kY�>:R�qT�����=F�p/�گ�=
�����L��mT�,0{I� zXM<�����/a�4�J�F�R�-�r�=����f E�]���B��^ګ��o]Ah��~�`Ğ�X(��VKj!h�?}vJ���C+���b5��n&���i�R��rԺ�8���ֱi�ˋ]E�=�)J����G��S�g����n�A .����ù	/��D�]]Ƴ\��\�e��J�7��Xz.~�h��t�Q�yV�Zd!���@>�T-�N��D_������	}�/�"ګM��ګ&�q%���`2�޽3B=oA�V7j�dh�S��
�f�oc	���P��6:4�0��^l�\�U焁�9{��1��`������t0]R�Yfx/8�Ƭt4��
��.�����4��$�|J~���1 ���U��Ql�)T�Q���u������M�f[�l���P6�6�hQ�"�)�"|�W�v�Ҵ��K�6�<����u0j�v���U1�MUH�R�-��Q�齎��S���&'?����/��-�D�O�5�����ض����U*Y�j�kM�Y"%����1�Kb�j22E�]X�Y��MyZ���:�+FG�P��ti�yՇcv��lw�Ys��`)mo��TP�Ds�؁[��)��D6���=��XU4����Y~�w_!mH׉,��4�ͼ>�ijBa��J�j�V�o�2�����¬�����-~ŀ�aB���0�-�l_�ۨv妰i�3���&{wE�C����Ե-��ۋq���|v���ы�3���>g�1~0 * ���K�\�{|?�N���g��2�I�o���Tfk�6�CuM2W��n�#�vu��.7�c\Z�j�I�6�V	q�O���Du:z+����D�~�"[E���/>uoy���>��78��0L��.�sjW��M��}�m����X^qp�>������B��@�"�1Af��ơ�,�1k�-��UՇLh{��+F�}����]yȤH,H;�꧹�O�Ι�h¢ٹ�HM�)6}��d#����m�)߇X�v����\��8�ŗ\au�Τx+�-��2����Q]0�ݹ��o���B�V&�$����'�wp�a���}�.���Y.N���a�,)ioԔ�1K�RNR���;�Ņ���0I3R�"�=z����!�\m�}l+��<��t����xv���L��X9%5�@7�ۗ�c��7}
�Qc��_�I�z;�4�}�~(c����s����~b�0
��dv�#\�����!�~���#���9�rH�g�d%T�m��S��{��	f,���W �QA�}�	S�dh��n�!Y�,�#jp��G�U+�C0Vڠ�4�8ͅs^�U�}�;�4���h_� L��=�8o p�Bh���m�q�.��)�Dv�|&� ����w-�Sr��U�j�GS���;R-�V�����v�G�y�ͽ��^j^W�|��W�w1^�pJ(�u�H��y-�XdHg� ��@�6��ʠ��R�Z�P�y� ��A�%�$�)�1��W3�m�t6?������f�F^���y~��+�:���`�^<gѓL&+F(��$��s�R�pK&Ǔ��P|?R�i�?���q��'�O�*x�_��A}8b�E���;�'�D.C�hM�������W3��[˖+I����6�)�y�5爀��w��#%�醒+"��c�T�8n��1|�u>U�e���d�&ZܸYvIR`h���R�X(�����U�-$b5,8\E�S(�ܮ�0O]
�i��1�+�5��Z�{;�l��?
I|�V��3ᵉ`�#_dr��4���X$ܦ��y$��X��-_�!F7w���i���j>t}�ib��ϲ� 5�rT��s�v7�u\�����I~��?kw��L9T��v"��m>��s���k�4ܩ���ק_�k�F<�0D��	�y_��b��G	�������V6Eހ�}���?�`��Fb��g4d��I�=�]� �r��4�u�b6��n�B�|tuC�J&��{?n���2��ڡ�D&��Qn��Q����- ��m�x2�l�J1\����̢Iِ�'��p[�B�v��
���zԏ�δ�2ѥ�d�.�~�����mx7��-�J����U�;���~b��B��������M���I�L�����M��p��`�\�;��s��榷���[8����KK�ĊG��
;��5H���_p���~�=���#
5�k������A�i��2 ��é=��.��}���4����olC6D�4���g7�θ�ƈ�q��gt��#�J`'N��E'����Ge����Kd��`��|'.�\\���N����^_��ğ�hꑩV|/�,o��!ǛZ/�>��YY��cT���,��n]�:*�����I�H�]E
w}o�y,�h�ťz���z5�A��}D������4)Q��RGhr����4�'��fC6حTt��q
-���V�1��{z��=3���ЙQ�X٭�z��V��N:D<{�'Aǟx�48f�oO^�z���3�QґŗʧV��2
�|Kt�TBGZ"V���b '����F���Z��Cw��ϫ -�A���x��u��Ǹ�������5���)@%��	[z��V5��{٤-?����"�3{�ka��������I�49�N���B�J&&���K�<���u�Ax�.qȻi�L����2�Tŝ!ײo�eF@�Z�x4����{�z�7نg�&�%>C����B�>O�d�YZ�i��>>>~�/�9'#i��^�_��يݝ]A�L-�g����<�4F����M�j$EF��D0J��!=g<�H�����+���cAGЭ��K�*�j�&�H��f(;�,\=�T�D�:r8ٰ`
�<����Ɵ�#�շ%3]��{&��,���]���pD�1�ߧr��2vx��UwLE��Z���~�=�Ʒ���	�;t5���t��ZM�J�\��%�}��DCVl�Ucw��A�e�����S���4��W���Zp襔�7w��Ah�2����$U�s@|4a?⻢XnHO�Ĝ��ZݐQ��n��˒1�"�{��X�P?be�;\���h)mL��$���ҾA����BʗS)_�eZU
Pi?� 2ՈI�F«BV��6���:L�~���ӊ�B�vI�d07���7��6Ehçe�X�zI�'�Gb�}�t��_"-w!�M7@F�1!��wD�+����xbm��Oo�����3�'�t� ��!�YY���!#N�;�<��D�� LW�w���P�k�"_Y2G5CӪX�p��J*ڟ�b<:ּ���F�0����5l����d2PaOxMs���J���Na�s�%�l��o�h��:�}nׯV��X%������y3�B�s�˷�71|��;;���.�{���!Rg���*�9P�齫����č����(����O"�^�K��(x?���UE$�kKPDz`�˛'���7n��N
Pǀ�e�:Xr�k�b����>��T� �4�э];Q����|��W{TT��T���m8�6e��U��vT	���q���!Y7��G-�<K�8_�\"�C?�
\�F ��3:��bف��"�0|3���oq�X&C���ӡ��A3�؊讎{WX��� �ܬ($|P��=�o9U�$�._���	I�8CP���q�Xc�DAL{~��.+K��-�".ϝl8�,��i������������ٚ�獐�Ub,�l�yV�S���^q�2�UZ�୍�EFH�sb�|��
P|���M=�G�Y�"4�����jg��68�:r�����ͩ�,}9�m�@���\�&��\��'��2�6�uÙK:C����CHژl���g<���UF�w��
3�/����
��ާD�I���r���ɢ5��6�g�"񯈴8�Nî��j�IID���ns�������S=G��Ԛ��pWx�� �� b�W�Rc_�����]���&S0q���M��k�e���������YL/����`�HU���_i@�l�z�^@���a�d��E?����K5:���[S���LDLDF e�=����K�C�����ǂY<Vˮ�C ���0�������P� ە���|g�����GpҶ7~5el���Zd��J��)�ŭ�}.F�t_m'P~c�I���<��Ξ_@��!0��$�!�B�^��Ԁ�h�	�9��㨞%6�TJ7D�4칵��@͡�X�ś�N�ڰ'v�
��k~�+ܥ/�P8�G7��O#��9`���N�.;j.�` �!�.*������� �1�1z�I�y�r:����r�o�@7��Ռ���P��9���N��Gk(���l��Qe[Ӏ�61H�Hvy��'N���z�er�U։/P���R�!n_4S�{Q|�w���Am�zzX���U���?� �}���Ռ���Xk�����w�7_bk�����?˧�d>���j�^`�\G��AJ�sq�l�rj
�����}���B4<�F�`������2�z��M_AWv���Ȏǉ_�\��r�=���N���KGd1�ѭ���-�9fBزa���F
���A����D;:��n_� Hc
���|�`�œ��MCIW	O���
�ty)�c����jÜ�32���NL0=f�� V��7�-(�l�!��Ϛ��'�[W���1��R�p�ht�t+�'���.�Gr8 �Ą���F^����a���_�����j�����d�*v.���"n��P�����I��]�lP����n��z��똶����]�L��(�G�uOJ���+���y*�O�ǹ�n�͊��Gu�4�]�@M}����9ATv��Lw�xx�䕦���K�߮Ѧ���q���N�e?=��#^�{ë}rK��dYƇ�����*�QS"����vP�0�ft�>7!�9[g�R)�_O�~�q�oy�)d�����4��mE��?S�o���cc�A���a���id���T�[QdِIO�|�(
w39�?�'V�ڣ�/�fK�G.�k�l�1�|�ź�;	O��,�m���L,��FW���A����ݑ$%{�+np���	5�ϫ���t$�e%:�3:��b�7�H\_G�?7w�Z�J$b	�h��u�|-Y	�����\#�}��i�����&�*]^�\:R�5�R~3�ry8��_��afo^�`3�E��1��&�jZRPK~2�s7Eψ�:Yk���Ԅ~!T�3·b���o'O�/�����L�m-�5}�M�E��	'��-	�4�L_����pA��� �kh*ή��cX
�7f�d]}�O��f�"��.��=�>Z�S�(��T��� �)��o�	jd;?�h$m�Xȣ���#�D>���R�3;J6wl����QOW�߁rC�b
��� �,.��-�A0�)B'c�%���Q��*��K0�^.�;��;6��Y�6D.�>�t�y�n��d�P�g��{/�Gl���?8"x��rU�7+zeZc�!8;��T��n��x���3���x�X���������4�Ś.M�G�Gayc/L=3��v��7���b�u��c�yH�Pi2"|��?��&D�|�/��h���V_%��1��1=	 ��/[�뚁q��J�gؾa�Ö����4\��&�!ɼE��آKA�#-ÏS�s�~��K��PL3Thj�5	e���4N�o���(,�W����6f��>�1dي�-,Z�mPES!��������8D���c��f���K��Lm �Ǡ�l�Ⴛ)ͥ���!�4���砣���Rm�x�wp�Y�WK�� 0�l9����bŖ����7��XlxVHYEB    fa00     cf0`�'<��� 0~_UU��i!Kl����Q�eN���87��F�������]�Ö�F�Q
�X��b�'_���4�/�Q9b���Y��Ʉ����A`ji�'��g�V������*��]jw^�%fP�٬��o�;��.���qS֩^]���]SVQ��F�5���vT~]������*�R��(\:���y���j�[ w�K�|�����kw���t*d�p�F�eaPo�h���EBg4.�['U�/5���iɱ�b��p �����X)v��ugN�T������`�iج�IsnI5��)��6oQ�4�I��w��]<1l�8�:�R�s{pN1��Nˤi�d�l��i���b�����(�s��s�46�����K����=����$ArM>��(W�ۂ��'@�H-��{K�esjz�aK�s��z�K�C, .����eH���a7$P:� ��m�c�`����*�Lh_��{��)���/Lx��?��>U�
5��q(��}2� 1M�j<�n�����_W`�GyV�؅(�Ͱ���1k��n[ǜ�Xpiέ>����с��T}��p�jE0X�;��X������Ic�	�������"I��5�q��(���΂��!L�Dm���X
}(�����;
�<Ԙ�2ep�FfCG�.�+�D9gE�*>�5��"B�cbO��N�Gӧ�eA�1~>��;OO�5�/?��D��2?��>��=�E�G��1*z��eLB�%�n ܆��K�{���y�ON�i����'���M(Q��5�.��h_!�����v�x-�Ja��K4\!_�l7�G1�:ʠv���d>�QOh����h�7�уX�H�&���v��1�m�{�G�i�:Lў�*M�����ؔ�SGG��Ć�ͳE?��p��Ъ�!Zj�O�솞��Bѱ�Ko"R�fW�6;�܁9�q��a�V$87׈�Ƹ^.��$��;j�Q���o@
�]��)8+%���qq6�ν����CH��˵;`�U�b\圃.R${V����{�l��	��~�~���v�؋$E"����Ms�)��!��ޭ�����y v��u�5�9(��ҹ�)��ޛ_1�>�Z�źNH�<r+|h���dP�]���?tQ�꿧���Z���^��X�'�NRd�[�`���@�<���?;&����S8P���0f��(���gS)+"�S��\ߙwH�!��1B�l/y\@8V���@�=��=������	�G2���NR��+�/��|�Ȑo�G,���U����Z
	&
�����DL�^�ʭ����˪�!��o)&����w$\3��-�c䚥��6h��wP��krFӚ;�MRW�e̖�S�l�9��؁���������I̤sJv*ǌYv�S)�h�wW��\8N0KT�����Z\M�J�L?á���E�-�W_�HN4}�G����$!	<��ӧI��x�<�4�+5�p'�]|�6��6��9zҀ.P��=�JbH�w�rf�~��|�L�����B�=9���6��յC*8Ʋ]���A
Ա@�;1����#�P8"c�ZN+�EE�����i4�WC�E� ��� �6_SM�u�%�{�Mt(gw�b(��~Z����g����7�:��7�M&�/�w�x���m���Uf���P���C:�XP����1���PL��n�U���ȝ~I�X�K-�H_]��C���O��#��z�<��S�=U�F�y8`�~������Z7КT]�&|!a��:�]��?��ܙ��9�䕉�-������t�U8^`�����E�[��9"E;�8���!�Ҙ���!�Ϋ$��gCy������7�Y¿� 	��wyCă0�ԕo2D������< �\D4:�+��������ӌ� 3$�e��{�R��4�JÌ�Y��w�X|P�^	l��	�Yjv	�N#({M�`^����Z=2�7��8�s�����#U~�����_C��TX׭��f#��4e���RuEO@�K�*k�h}�TF��yvka�=%�	�˻`�X^ƕ�UF�HB�(8�(�VE��AQ��0�=�ε���u����ȃlg7��q�}i�bP�{j�Z!ڤ�"m�������K�D��o��r�~�������5w�oz��3Ԅ��cZ� <��Y�ʣ(��0�����"3�5�>�`z�E�
(1�ڴ��Q�I�f���	97�E#X�T��]5E	�F[�j���1�!�8�{0:o2H�͚�z��V\��]�&c��z[;z�[�W>���ѭz���މ�*�КƩ��%�˼:�j�{h�˸��
�I��iE#/�1~��-��Fu�t�`����L��K(�{�������/��K�B�a���8� �m�5*�� �_�d�$zV��p�e��@OJ�Z:gO�[a]X\�p*��#@��@�`�jA}_��H�9a��� �	m
aP��ڲ�H��Cez�yD�v��}��=��t�X��~f�ȿk�\6��A6�_�[`B��t�[�s�Dqu�Ҳc	��ÕO[i�	іz$�Gx��f�K���� ����cָ����wn"��/,�ua8N��BY�گv��uy���2ba��g	PJ�� �"?�Z�HC W�#�?1��aE��
��&��گ�������_!���pR�|��L�8������H1�g�8�ޜ���� J���Ѽ|�d���y�aޯ�9A�V���DM�'<���u��Y��i\<rcfĦ$������zUwJ��_��*c�0�bL�-k.�K�z�P蠳̾��[�9Yg�Ê��Q�0\��i��w�yl�ZR+���]��?�0���1eww7�ޞ)=gT��Qw�Z�A�K��$��73Ds��+)��� CS.z�װ6�~c>�����o�$Qór���D�bZj���>��)J1
ԭ�c_]錦|�꛶imS7�⬨�O���Ѱ�?J��m��{5�xȉ$g��������.ٝ砪6��{�|�J��<:z�-g���#8���k� hQňyX�A�����S2��[:�"E@������H	���e�sm�Ŀc��� �6�{����ϙ���� � �i>�C�KG�ƿ!�l�l[EŏFv�e�-0��T~�&j���}�6�[��$/�! �P;<�Ö��� ��▄&}����P;4���-�q�ڐ�d�|�i�(ԺyB���a�� �ylX3un�M$@"��wR`�XlxVHYEB    3981     4d0�!�~]��2����9��;X�n��ذG�N��K|�Pg��.~��O!u�V[�f����y0,z���i��^N�Y##�T&�#?�4��2l�����d�n�'6�<ٖB���:�j����}��"�(��yn���e��V�u �(ZP�>�BHO�+�iw-y��*q�8��*.x�G�̦�ӕg�o/C� ���Ѝ6�h�i�nkV�u��v�b�x^����FGZ�[Oi��gn:�!㣻K9��/�mhI���������%���T��6n~�}2���iZ��`�_\=	+�u�_��ue:_�!-䁽�=�j&��S�yW6��G�lq�N�g�%]Q��^�+���.gt0���4�*%Ĳx����j��$��aS!��yTΞ��y5�q�r;���)!/��vbTqL��{䝿ʰKa����Zq�e�MI<Bb�0J���� H��Ü��YN���W��ch$,[�gj�����.�fʲ���Z �h�+
jRd;����ɀ"������w�Dg���m�i��o^hLc;r���q2������S����;Z�8�]����'��{/#��	
ѻ&�Qea��<dL�<���,����6B���\�����F���کCl�L��W�ؑv}j�~��v�5	Ɂ�P6G�9	���B�u��aU�M.CB��},aL��@'S�'��z����L��wn��C�-�N�V���-}�v��B���c-�@6+��(�P?�����T�Ո.=�T�!�A|~ݓ��>�lU�`5�.�9�e�յT�>��fF����"��oq�A��n�P֩ iao�ޤ�����(<ǴB��^n}�ڪn��I���bx��ъ��IL\��`V�'��Јɋ}���"L*�脠c�!�P\փ�̀DÿrK�R���{�Ҡ>)j�a��=�l�&��P���at��������=���YD�dO���29�o�є@�מ�dQ�؄Ű�q}-WϹ�/H�r�m��Q���d��?���vg{*�y��p:�Z���d��^ۜ���gꢘ���nxE�P�>�=�$�4���2�Z����B���#��e �cr�o��'�b�d��~� ������Q:��/JM&U]�C����۷���c3�&��_���'J�w�@�|�[�M�M��yC�>�[�g>eq/*Ƀ�h�P,�Q�