XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���).L<,�G���jJ�D��vX�@!���|m���m��@��t�C������#�һ$���>�|�b��;j���?��.S �o��q`E��/���t�<@+�a/�9����̣�CZ���e�.�� Ɗ>2�+����ᆤ���k%����g�p{�|����;Ya8<�Hu��;�'l6�0��a6
G��@�w��"�9g*c�b<0\��.I����v����� �= )�hI�X�a�R=2���~g���B������^���Ā�ε�>S*���'rk��1𡇬���y�8`se*��e��v#��5�Bu��x3�A�Ġ�S0ܛ���a�"������2�wN��_�5��	:���8�.���H�����&BÉ��Y[w�2��c坕M]�
h��Ǖ3ps2R��l�P�P����ׇ��-Q�^�����hJ��}�����*�3��8^�@���5M�·�	�Єn��p�X�_+1���i��)�^'�à��G��[oU�&$G���kh�P~�>��%㥦ah?+SW<?ه��xxy���٦��V��t�{R{Iy���{�{|�;��K��Qyh�����L�Ɲ�X�ىl�ruÂ��9Ebl�4P��8�K}�ц��p+9ڷ����9���Z#[�-r�^�u�o��� �}p@���5CK������K�0�RD�B�tkP�=%~ ˠ��R¼�?�|�fDP܌ج�y�؜�A�W�XlxVHYEB    1641     860 36���p���h�@~|��lm�����ݳ��/c��4�0�DN�~D�nXf��b��m��
(�U��V�+}dd��4���P�N�Қ�y���9CV-[��������7]�\�6^
y�ڵn+���J���VP�&{l"3����x��I�{+��9�M^��G'*U��+�A&��2�I����VljT�l�[��l&4@�7G��,3���؃aꑅ�p��rBp���02|r��t���]rK��'@�"A����q��y5oM>��	%mu�!���XO�>$�*��m����e}���ؗ��:P|�����=��G� �ǂm"���)��F���&Z��gE�?�w{qL&T�U�]U�F����P�g;ғ��~��1�)� o�?5
��]����œ(?ZV7ؒ��m�_峚[%�)�Zo0�1(1�r,��ҒՋΐ�������X������=�z���q����}
��Hm���{1��;����x�����6ħ������^�þ�^T�ۯ�	b�wV�KbA���o[��M�y�Cu�2������ٽ��NU���}����_���4:�|���n̯U�od$�����%Ֆ�m�rb�=�P�6q1X�'8�(55ÑJ�����ٮ���Grʁ����%�Gx�vG�jBQSc
F��k3�kM�v��#�7O����鑌� v��x0���R0�!�_W�(W��X�O��s�ډR��v�#in�{M����b,k9@�뫾F��X��F�
I��|��8���f��]3F���k�m�1�h�##�U
�eձj<�F��Pu|@
z�`	MH^5WR��CPt0�.6+ɑ��S��y��]�?EwC����=F@���z��E��q7Lu�A)v�*���7��4����i֧��Dah�V�[��:���R�}���JH�a\���;*f��a���Ã�XGTe��[ñL2GG��Z��o/�� 뒽��*��)��IF����;(U�׫L|��]A�[�w/��tlO��Jd�`;ԓ��)Z�Wa/�Ź�{�
�R$6,�b��p[�v=Y�7^��Ol�|����W�h_��ț���Ht�*x��e��(��!L4:��-
/J륺iI��9u��*\su��Y���c���&��}�Jv�C����.�,�$NDk;��Z��
2��0�9+��-3WE}A���[�<�� �2b�m� tQ�=j :��	�./����AI��6��Ar�m���ʉ�h$����MQ��h���_�%m��+�u��^"@�qF`�(�e�e��rm�¢�d=���5\���J�~i�1�V=lT�������g�4Z�Y*�=�:��(qVBk�������5 G}����{3[�r��E���N�'�V
=&������Y�HR����7�t��� R����T��_�a�'��4\u�e��|����qW������O�1nf,d�E-T��7o��)X{��I��V�u%{��[sfl�<��YC�:oo�h�����})��z��X��%|3s�P7�����MJ�(�ҍ�(�O-D���|R �+1��̣�2x^i+ÁD�\Jo�Qg�X�>S�����̾�Z�ڸ�k8!��7g�Uz��RR�+́�� R�g�T�52Ŏ��{g�a�⪀��$T<Т�D���ѹJ	�l?0�n$ٲ���+������X�lQ~.�0%4�ǧ�`�~��� �KU�hY��b��4�T�?ˁ���X�C'@6z|ìp[�V���X�^;�%��{�;�O�#�|�7�����#㯂ኴ��H��c\Z�n �	����\�=r�F�s2�؛#&/%f8nˏ<b	�s��Y~T�|&�:�'De��{�T}D́!gs�k|Ž��۔��G��C�kc?pTV,�����b��N�V��M����o����$ܕ�-��Wi�o5���ڕ�E�َ6it���T�i���.�_�_*<`�
��L�Q�]����L�M����Z��ԣ�����3DZ����Q��$:q��@6��(Y,-�°�)�����c��;��C�x��%YI@��O�B�χ�f3��F�4N�T��p