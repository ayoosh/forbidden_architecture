XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������1m[�j��*Vp^� '	0Ov�k8i-c� $����@Q������B���Tz�>b��n���<�I���KP<j�mjIuM#C�0ޛW�l 6X)��V�u%��hN]�%����q8����Z�;^��5Xn�!�ق�m�;��F��l�K◢�y��4����h����D��~3���\����W$'�����&���8@��n��>���N1�mÂ��!KOv�p�Ӓ갳D��'*Kl��ZP��w�������G����c�m��S���m��*���r��A�zK�N��G����.�=��&̤�m�����*�&�(]�l�FM��:�ĭ��d�^��v*��"Vc��
V��rO�]�lI#Br$n[�) �U�����k9y���T���1=
��p��`T6�R��c6V�C�M[S)B��*��������ΩV��.��;����ϴ�����0��f�O�(;�����?H�Lv��i4��r譹
+�K}�!0�B5�>V�%������sӲ�g����a>�������:�7��=��9$�޸i<Qd�%2������u(��7;��t�7`��Ɠ�I�߾��j�]<�Zr~����AZ-Tw�dP���������3l�z����]О�f`���Nw?�Q~�v9�Zd[>j�@&���N\2V�:܂�I5�
�f8���ލ���\s|`��\	3Gh��
`�eQq�c���1�
�$W�ʣ��4�XlxVHYEB    fa00    2220 ]�w��菽��I�>�VN3cǘ}��>G{��>W��.���2�r��F�['솚Ƨ�V�"���-w�R��^0�B|����|�ot������!�w'B�ot���@Q
��:�'�փ${$"�HAJ*�~dtZh{8����G��t#98�����n:]�y�5��:u F���ŖMM�n���P��7��(2V*U�[OI�G]	N�S��G�l�꿸��U3Lڦ�1j���8d�l7���㲂�9ֽ���PnT-�i͑�d���߿�� E�M	�#$��@b�����h�Y��z�8[z4@�$���գu�l�o�^�b���n	H�(fV��uީ+���l��|�j�a��L��C�	�$^��!�nu�*���5��iD3����*y�49k4 ��UY��Ya=".�2������K��Ab�>�~�T���m���s�sON�6A[t�m�
A��'9��}�����닼�I��~�䠷�(.�.7&���s����϶Y�Q����-�pvup\�?1���;��=x�@�f�)5��]U�d����j?9��i�{�{%���r��&(L7���t�Ǭ��!����W
ek#���s�@_�[�4rV���p��=����x���Y��V�A
����:��F����N v���2[���;N<^���"���^$�ԛfB��r�Q%V_�E�ⷅ���X���M"�T&'o��WI#�QI���إ�q�������I��BU��-����p�tmv��7J��W��lXB}�
\+��5em�ooȎ��͝d%$�����&|v6��<�4Cu�\'0<�,��Y�e�F�܇�����x�Cq ��:(aS��Ҩ)w������d�@4���O��*�x�^���|��kMMszҤ��\�.��� R%���N�#\ή��n��"��*�0 0F�e�����gk;�,؋ 궴w�@ec2߃.�$y�0T�= �@�\�>�]+���]�^�Z�o����	l=^��H��Zc]��f��@���?�q[�[�5�~F� �4<��8c�Vq���-Qw_]��6߯���3������$�u��"}�s�i�(L�i��f3T�,��6�O{iЧ�~�p(Y���R�tĨL��%�ng�p��@s :7�G�bP� ���A�:�M婝�GZ�rh��J�+4�"�!w2ȱL�cc>oXF��'})���	���aQ7��CUIq�)��={Æ~b8U�2�[�qJ�E]~�5��<��z�{IoK�&�/�������������6/���}��{����y���43Z��k�����S��+]���.�ᝎ�_�w��{�=����`~��������b��V�h��?1���K��wE����.�N_N�Ж�6������
���l��Ӷ3��g�4)�����_�=�R2|?��z��6�l8 ��$/|}r�;�6`pդ2�];f���pVB��Y���@�Pq�؊V��g~ܰ�V]���n�eE�=�#�Y��kWm�up��'%g�-��-]�o��~hRj
��2eҶ8^eϪ"x���l��H�gU=r���Q��<K�@Oٞd�Wɿ4��;6�����H"5,�v'�j�uT�u�>��L�8�r�rC�mS���2��G&c�%=OdTG�pWl�v��×�.�hk4ӳP� ]��ef�p>6\3g��O ��e]�P�-ѵTX$��ALx�V�P���/�����Llf������-2 e��L�!d>���#f���I���n��Ԑc���0�ǌ��6����e;�6L�I��)է+��t5����2�D�i��\^�J��eM�"'��B���ӑ*�f!�E h��9��[	Hج���R[��Kt�&���W�)?�g��c<��o'd��8�&ȶ�
�����GP����V~S�!Yw�]�����4@���0p�S��xI��p}"�3P�S��Os�7OTϲ� -��NU=H�R�4H��Z��Rv��o�BuP%A���׊�[��������I:�lS9&��q��!<W��A*���]�gR0����Ҷo�'��M����T�K�M}	��e������;||����|�CەM�	׿��8�i��F�C���(>�&�l�~�̪Imr�U�e��
�B��j)�{b�tΛvЀ�lz��e��wU��������圆��\�'Y�B+*�0����j,a.��3$�׊G�v�T3�]����ߨp���吥�aVuٍd�R�c�]��.�|M�a=<;>����>��3�sɎ�qԍ�'�>� ���|e��q'g��r�����a���GG�_T�j�b�%�8h��8��;O�(�C��Y�jK���{΄D�%�
��X��}�@K�%M�C�fqvX�H҆7υ=�+�H�3��{�r�w"^�G�CÞb0�9R���#X�Y�W&�<^>�%�7��#>������h<��K�NN�"��_Y��!�d����p�0=R܆����>�!y�U��nV��%�4�i/KQ"7H�H��A��X����v�|f����Y�T������щ~��.78MU;p��8��
��Bu�'^���t�8ZڤO�ă�wd9��g��ʱ����9hTt}�+���ȵˍ�=�%��7wW���Uؓ� �ΐ�T�݋�+2&���I�@V����#CP���H����N����&)>��1�� ���01�5�I�$�Z�/���=e��d�RÔV��ڛ (���)&>�!`�/�䛓+�� ��n�&$���2���w#~2��ܸ�R��r�e��]�fE/��e�9��ﴱb� �?�I7lM:��$}4�!}5,9,xpq#|r�"�݄^��)����4��`�Y�%�����ɓ���>��̯�Oj���vE�����W�hso�G���pg%F��%W�Н��Ng!�}c�ܸ��lf�f�\:K��� �V�T��	ɾ�D�.���*D��y/s�n�]zD,�@�����f^r�D&8ԿL;��� ��L�����ȍ��2<R�o�V��5�~�D<�Х�j��;k{���땕Ӫ��!��iY̘���Dhcdf��z�_��[G��10*h�ݵ���%�U �ػp�ED'���@��x���'�c�:�!��z��O�f�5���+���F�H�a��^��}�J��b��Ӎ@sȈF�H�_�2`�n���-��J#���u&�>Fu���[v���D�0y�x�\4�z#�o��ؚ������x�H8ԅ{s�}�K겆q��	�o��9^u M�z/�����&��).� ���-}���[I�`+�W]��� ]Dl�����J��${}o��:<�RrRW\�Tj� ���<'$q0창4F�x}>�]E���ԧ��Ê��Y�ovpd2��#���JS9eXU։%��+ѱ�BP:��M�~#>�f�)�l�D�����koS\ڑ������l��w�$C��yۦ��P�[Z�k(��>(�*o�!J~��R���T4�#X�Ӯ���:��)]}�����iۧ���x��L��PvI�/�E�x�@�x �曟�����+k��@O���gMrh��y�����&�g�U��G��T�[�o�U���_W�0Ў3�D���4g$��
�A���ua��ݍM�V���}���}���W�D�oo�d�m���B,�[=���	ܔ:��qnp�p�%�ŕ,�M�[���W�<�	9z!;F����wIb��6�fo�/��>]"�vZR�:_�C�x��?�x�����}q�	R��T^�MvR�鮡��%�yŔ�ϳ��䟀�����]����xL�Y��hqFf�̥�|�;�
<NE��]��������!z���U��OY��������A;߷��LMb�ϸA��4Z?�躿�{���:����p��9�c�g��֙�N�v�1K(���� �Q�*j^D�-e*T���5d{P��A�I���rIx����|q5�F��9��@��<��[@Y��v��r
n�HL�R������-Bl�~Ǡ��i�(ބ�!�����!�>�h �N�iL�g�}�c]a�ݘC�D6�77c����osī|e�����@*0��Zn|�m� �p ������UyO�OUt���eÎ��+�кz`�{�@Wg�6פڕ	���f�^�h;����%�k>K80o��H��Q�Ӷ�A%^"��b8�G��5����7��.p�Kd�%^��=��7L�����>3�a2V�sn�����! ZQ&	��0�f�36,tn%{�o>]ڼkC��k}���x�S�0H�ུ���R�<�u�<�<�8��	��������gY�����y����\��>ʹ���GXF�5�)GC�R3�_a>�@:W=����V�?
fΙ��S�t��;�:�Ϩ�b>�~Ĳq���E/N�%L�e2d��d��<��i38�+=p93O	ll]+��m�w:Յg�H�Ɩ�q����B��zx��v3DMJ��y+G�S�8J����]1f�Jv eE� �T7O��@���@��a̯ٸޢ�5���C���3���ţ�j��;��ͯL�:�);��?�d�y�����UD��Ex���������1��
��O}�M�ɡ�Iܸ�ʽ���A"���"Q/O��g��h���F����l7�x5�Δ#�&��w�]��CTMKD;��=���̄H [�rw�_t���c�yb ���H��q���ug�V��x���1�~�:G��Pi.�B��x���`�l��̇��(������gn�V���.]�q�tm���u�����	g'�b��@3�O6��g���y��m�*")��8_���[�@�>��L���dA��M�,��a;F����3P���)8� �˔spr��m2Ҽѝ+֮���l�9*�0sc͊|`�ܭ]TH:vP�����>?(����z=zk�E|!�7&\d���nt@�0���:�9�sY�8��	j��bו���|+Ny����s�t�
x�aQ���EzԤ��ɧ@�,^�>�V��9g#L�ӟ�F��)��������n|�.���rb����}ϖ!���(�{����ԧ�������3����obpc�	�S�4e�k  ��6Y��L%FEG'9�Teoөh��}�!��Ż�}ZR��gi�Ss`�wA��Y�@�]\�I�� ��İ8�ɒ@�ݘ�W����>L*\�$�������ݐ��N�t�噽�<��5hO`(	����w��ZHtF�JPu=�������SR ,;�5��p���ڤ�xu��1�t���t�U�\���:X��1�Z��M!8����$�l?��`vAD���O�������%+b}$.�j�u`Fk�9�<������6D���a�i���a��{dEo����l�K�64$�Y��Ir��=�\���>��>��}$��J�X �_�[�$q���o0��t۴��f���y�v��ʭ�,$/e�.6o��.9p~�4�ۢ ;���)@\VY�ZR��P����H�*����s�ԟJK�>)2����X���:.��s.m�2�U�!9�J�ŝ;��a��Zu��`�p=��~���JW>�9F�Ҿ�~$���d���2X++}���=�5,���)�2�Fg2{�a���c��&��_��Y�l>����q�	5#����w�v�:��� ���,?��9�ШXf`�E���@-qb���ĭ�['�9U⁹�Ή2c>"��2�.���A�}��1l0g�T��,��!g;�z�i��`����W�bq!��a
�`�!�K��N2w��g������a�3m�ͦ�N����Azp@Q^��⾜�_�F݊�\q	��MԽ�/�y0*����'bl�c����)���p9���>����g���7��g2�?�k�T�a*�8Z48��λ��=�9O%�	�Ti����M�~Ӫ4I����c
�[hv�"�<��V�8���7AkՒ���u�����$��~侞XYxA��q�^�����7<	�b�k�Ȍ������M���N�Ȥ�m��N�-� ����َ������9�v�,��)�����Jԣ�U�]W��q��,��^���@�f�k������+^߮��/��A�ڧPڃ�3��)��N�_�\��;5��8�L:ˆ�Y,O���|��cQ4��HƴރaV�P}��m��ZE��߿T�����1t�xA��Aϕ�Hn&����^1+�7��L��y����B:dqK�^�[f�C�W.N�pA���|r����U��M��bǗΐ����qǢ�����&��Z�:�_Ly���j����K��<����8p��8��F��	�_�Iƈ��C�idA��0<�/����`%01�t������R��.�B����4�]H1(��8�'S�?GM a̜�Y0��Y%�,��'9v}�?�� ��f�/b08"Q��)G-�ePXw#q"��J��l�[����֏��E����N�3D��_��L�,)���7��F:��n����8�ny��XE")@�H�����2�~��ꉛ{+�)����E�����y���d��$�'��	Gk�N���]9��x���A�.��Q��%�%����B;����|�JC����!0.�7|����?�|�l��6�al.9]v��x���	nyhdeu;��Х�a|�6�Te�T��k �gM��ӻ�,��5gdz+%�&a5Õ޸D��%�I�嚧�����"���K�BMv��L���p�x)�U�	ŷ���>���+_�0����B�'�n��\���jj]��Sc(��vc�E�nű�>˥o���I�#x�Q|;�Y������U�&oϷl��ݡ��>n��^f-�2�`j}�0��VhIG�.C,~�8�>�n��yHI�8f�m�4��u�I�+���4p��Z����[.��)ox��ߠ0:6X��wޅ��Jk4�0t@���I��؁�7<\�5մ+k����0���R������������K�\m���Q�EWo�ZY��c]���CV�U\��&�N}�������}�w�c��j�y�k귨{���2;�MC����y-tm�%��c?0�[EPd�Rwz���7�oS�	��r���xf�f@��ir�rF�5r�Z �^�S(���j^ⰡH�!hg*��RNZ�gH?aa��T��H�����0y"��bC-������O�4�ʅ�4h��
l��?�wjL��mK��!�� �M3�R�c��.������Ѕr)2q��wAJ&Q?E�$?Jb;�{�l��Mo��'��~q]L�V�)��#q�Nv�T�)��9j����u-i�T�(J���HI�V���͈-���iTH�m��8?�Z��p�4���$l����$a�_�z��=���6G�b��D���k�a��[���6�zz7�L�`�}���ބZ��dS.�!���qL��0;Tw~S$��5'}�,(cR`o{&�n3����q���3�6(��S��OK�f�Y�/
����᛽C�P���&eP_�%vK�\��ױ��x��B��8�Hy�zr���o��D���r��]�m\���V)��<�~WG�u��q&ooϞ�o_~�{�}PZ�2^���?;�)��4�5���OC�?�^M�+߭`i�����@�}  8�8=8�<���dd^u��E"�f�\�ƒ��$g��/�C��Y ��x��LQ2'�kr�H��P۶ߪn�%�'��:'����oj
���T��,FB���e �}����p�������N�I�W1�$�&��30�&�Yใ^�Ƣ���U�|J!+(&@�'8 �X�g>�����/B���a�pa��RK�������D(�²u;�Y�����u�*'Y���r}��&՜��I�{i���^�Jmpq{�hOyc��ts�A��i�(��1s�_j�<���!�,w�������|TOD��{��[�#�efN��6�~%��B�S��͇O�����!���t끥E��_a�`Ĝ�,h��*@f��x�;�J�ň��[������|Zf5k�E���c����M,��l�>�g�z���\�F��3���ڍ�؞*~�T��]�����0��][���O����F�d�k�Ec9F(C���8'Ɨ�搤�\ )�fdGً�QӘ_��%����J(��@���S
��N��-���p>��������^_�vA�,[~�#��H$'����	��C�!�=���j�~����f�\Q^�}��A��JB�>�　2��/)�>��wl�#ϟ4܈�ɍ�<K����[��B=wR�����E���D���g���O���'(�������z�`�ӥV��a5���Ŧ�ڞ�+�X���Dݗ�)qv��6/�� //�^��x.?��?��%��{u�m�#�9�#���&0��q.���z~�Z.(;[_к�֭�ꔳ.8�.(��FXlxVHYEB    65f4     5e0�w����r�������R��J���^�$��A=�2����5�u��D)]����r�֣��&�T��\e�g��w�����薴n�uA��>X�HN�v�2�s�[c�F��D'���0��9)�r���i>���CV�<ã?�B ��: ���E�e����d�+�� �F�G���r�׆kM㔈U
�&���wȧ�6jIS� Qrmx�0��%uT����D�z"E2��ͪ�xꋍN����8
v�k/�� b���g�7�;�K*���5���Z}>��p���O�pC�.�x��l5��(��`
d���c��KaN�'�&q�z{Jڌ�.��d�g�dq?�XMר-2#�glr����3�҂���>�q�Y����9�=3�ە�e��)ЬG|�n>��;�0�qh�Ǆ�Ϙ���Z]��&�3��qn��C�X5@̀d�:���G�>��~_��˱{���=�d� ��L' Z��!���:��V9��z"|�b���v��Ȟ�22]�&9S�ʡ��~a�Lwg�m5�ѥ�l�׳8�f̥�x3.�x�6�,&��2��O6a{��XUW�y.yTz%l?�͈�">C�TB(�ږ|���� ��ˏ����_7j��-<�!�`h#�R�L����PT�	��f:�,�tz�ȯL����Q��!E]7�<�@ŕ�@�fg.}�P���	1�U�}�����5�_<��KU��hM�|�����(gq�[F�)��n�3wWLޚ��6�fX��~ 	vL�b���Ց��ϼ�o[v�:�b|Цx8Z%д5�/�CS^3��W+�	6���ec�j��A�=�rWJ^^��S�\�l��k��s��W�eκ���`���N��(;?��'�U[5C1<�|�X�#���F[DI��`_R��'��=Ou�����^}��Q�yܼ�
��ש>����46��h�l�q�I�X��/T�"Q$W��=��0n�p{��G�����b��&����KR�͍�@�˓g8t���@��sܾ\�x°��3#�W��2�̘n׃�(�{`o���M�ma��z�B使�Ty���2$�OԨ2h��.p����v\1TQ��]�* u�����x��Ʈ���G��&Ǵԟ�nO`�An:��l�z��G���En�N8u]ʚ����[�Kj��*e��X��0���`��A�4L���� }8�$�{幻�_������߷�Y��"j2͍\U�MO9�|����ӊ�QK�PO�Ei���=���������$�)�&�	��qx��U��'�B�_��_�CS�pӈO
O;:�����C�V
�&����X���6����;X��i7t��7OB�6l�v'���Boά��NSP��_�B���{#�;��@�3���1���:�"�Epe�O��:�I�v4���].C��L%��_<b�n�����.'>��`����]�o���\��;0�