XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�NZ�th������XM1~m�(�	<Ī�9���r�D���^�	,{�mפAjK���$}�V�[�jy��,*-mJ������}M�]��<2��}��y3KQ�'�����bkc��
��9�ɌG�!;���H}<���V($4�b�4�N���P���(����W	���̀�fk�%@�'5��*Y�ZJ+r-UK��e&A5|���OtF��"�����T�`�;�@Y��x̟����Z|>6?�������40��t��xU0X~!�����e�fs�$����{��)��Ѿ=f�e4�a��B�B6�K�I�m�0��������V�x��dI��/�Ez{�SD�,@P�C�>�>p�x! C���O�YD�^M3�1[�LB94|���<�D�0u��(c8�Xvt�����E�)�ii�m�w��f?��!��i�J�޶<ol5a�����a^�u�.z��u��e�'�����d>ΰH��<�P}��_~��P�ؓ�%+�~�5@Z��T�v!�F5qKȨK#�5'jm��'�$����*����8W6��\��B�d�8�?��Օ��^LM����nwn2 i�9ܝ�)0r��mW��u��,(
Ɯ^���=]� 7�B�˝@��D!�3��!Pt�c�!<i����I�a�0�u�NPH}������뗗���3l�@��YR�w�U �섪1#$W` -�Uƚ���N�d�r&����1�zQ��*��A�����dI㞏����V<�fXlxVHYEB    fa00    2500\��gE�>m���C�gi��������=0@����Q��Kp*�wT��<����ͺ֏2BY�4�Y�Q��_,��*����:wۡ�y��eL�����pO��(껈j6��`L�q@�����V�	y0Q���SGRt���04ۏ�M��CSxa����=��|��n�~:K~~|Ga"#ylQ��%7(��OL����NճG'��:��a`m/��R��
[^�i�]�,^�~�Rp"gDb��e����7�\ ����(洢*�!f��F�4zr�z� ca�,����4� �߂V�;r�Ʃ��5=,��ą�E����lv�DwЍ%Ra�ڂ)�3�܃��sӘ�4d��IA9����g�o�z��������d������BҎh"z�k�m�V�j^�?ueKzL�vRd��%�&�K�3^�I����T�x�-�8�%Y�n�(�JA-����m	ec���Ⓒ��v}^�������l�fT�ѫ<��[�**�fLgN� �G����J �ME�t���|��K��AWA�)�j�Ux�Z�c�)Qm5�>�l��_��`:Hk��4-wl���e{���AY��� ����x*D�h���-�K	0׆��(��O�4�N�~�  :��l_=��5�"t�W�jS7�T��(�dͱa���
���O� ٫�7����髿tݜrI��Q����P��'棲(!�Ӣ�}���X`.�q��*Қl�	Q�X��TR'1��Ĉ��4���d�B�U0RDxU>����%�ճ�𜢛gጢQ,��@-�k*h���ư��62�*�+��'u�R$�)��sn�<�6P1���ӽ��'�l�r�(q{�{��>&�w�8�I�>m��]MoVi%6�����4��!��8Xُ��WQ&�^�wNT��zBP q���CM���Bg�&�aOA}p#�Gް>Uu�)� m���:W����yr.��'G21>uY	>z�����p��v�6�8`<�Xsu���8�Ε^+4�س^���&�4XE������l�Ƞ�^��k��h+����J�������4�K۴�S����@*�$'��:�HA��#���2�;�~����*B���g*/�3� �,��<���hYq o���!|�M��:��K,��a�;s[2ĤkKȸ*G
�.T���;{Ԯ�U\�-���['�N������t��?>
�ӑ�=U����eE�)qĠ���J%Qz~�"�Ά�j�Gn\�	��^s0�㼿��>��[ek�1Ԏz�� !H��&��l9!j~ڸ<��'`�9��:C�g�$�!a�|�ύ'�(JH�x��i}�d��N4Y4���2tҵ�܉����v`+�8/k5��J��w����z��x��{x�>��=->)i��A^~��Ѕc����[�X�4����_��͛W�@��<���j�*��PQ��D9� a�۟�cR7b�B��Ĩd���U@�$Î�񽾂�*T[E��-��WI@[aDH��1{v�P^X�1W��A�j}=���?l�Ό�A+�����l0�5��L;[���ĕ6�)�4�k�	��CF#���'�����qx�rbN�Qr�|�m%�hdl�uoҟ �4"�t�:���M�GF��2�At�9T��jD40�8��
8��d����-�h�zC���|T�qyM�
��kϑ�Ʃ��ʷmd�
�q�����B�GoQ"Ё�j�?�OU"8�)oRH�*⸓�dS�=K2׹�{@�%g���ܯ9�q/׶!���FA05��l��/	q�7��S�t�m��OSh�By�r���ݒ5+����&dn@�mC�f�A�ZG�xH�ff43 2S��j�����_��'����P{�XW�QW�����y��fW��$�b	�'�#�y
�E���0i���9�I_�ZKa�f��m�{7QA���di�~�v:��UJ�#�.Z�	:�h��Qt/f�/�TkN���!A^���jVpT�D�;F �/����!���o4 ��0���$e+����r�|�ף@�G@ò�@��� xG@ � �Vg�%�Q>��G�ι�~���Z��ף��[g9Tp$�%B�w<��C<��2@.S�w��0��0o���D��]V���KpĒG�T崉��.�e=�_�?��t��<j$O��Fb�;�-�a܅la��8ñ��$�����@�izc��gf�T��$ fA��w]Bjtۣ��'���]��PL�/�	���G�`ޜt6$P��~�_��&Ilr��!|_�|yR�R�ٮ����UpnMp���� D��:����YF� Y�������H�[���Q]�m{&��sd�)#[v�J$˼�n��/M1�>�u��t&K�:��kŗ�7�La��s�!�D���/g�5#��I]�9��u9�K���,��y�� �h���0`B��(��ġpPѯ,�2֘w�XEYD� 2`���>��?��k�d��<{-�WǤ��M>&_��&s:�'ߡe���)q<O��0���4F�4Oe��@����L"@ ��(E������߲�1��B�!N��a�Lw� �;u��AWxx�.��ql~�N�h�ǃ.gj8e.�����K���y>Bn����6#������=rO��������Vn��^,i;=�=2��$�#�޾QXh_�UA�"���
SA�Ĝj��_�zL��p`Kt��Ҝ�$8��]N��������D%�]�J���)׾�D��B��1�����E�_�[��"T#���r?7�ƼB��;�U�:�����ۈ��Te%���,o�����<:�l���H��n��N@���y`�o��?�;�4���o�N>�=G/����R5��W������)SQy_���⮷�6	��5�����e�fas��8���	��\KT۽]����	�w�j�\��eOS��(�\�1s�!�v3��Qo.I�g�%��Z�:*A�)[�c���)$����3��Ӡ"'�|��#&���C���k�"�����'j%{�>1ʌA��\kk0��?�W"�,��mKM}�41a2�>�����Sk��r?�`���=�4<��K1��l���U֘޵��W��>;6�3�Y����	�[fO!��.�Q��Nm]�<�+L� �r^�F����Z�3��r�P�h�W����0y	*W�dM��� &~T�Z�VP�>l)1!��Q%:�"H�<g�����������[0��[���
i�k���%�C��1���<258x��|�����"�qA.D�g��p<Y�YB��3UĔ��v�WΖz�P�O�6M<=����5��)�'Aʾc��i�)��K-��g|��>���vt���bT��e��%̢y���Y���*y6�W*�E(��!�H��NƨΚ����%��2����}��+�)i�a>�F���w��� �����l 8��)����V�5������T����s� l���մf9<�-�/	�ۊ��+=�!��__�o�7öq��N���!��LS������	� kf�A��f�v�,��L1�Ov�b�W�̻�h�)��8}��(��=ä�-	�*�lz�V��`�����Tr�:�����)Q��M�N��Z��e�_�1�ab]����-#�	P�$�{�~��Sz �&Oe���?��)T�#F�g�]h1��56�DB�@�!y��>���裄8eu�	�!�uz����I�����|�X�z�%U$Q:���>"i�����=]>�� 1����� ,K`���2���=�������sf�J����Us�-m-�2�oH�������׈N�#V��W`�`�K3e�"P+8_���Kk�?��C<'���q$��T���>;ǈ�!B�__�����Rd��^7������xt�Wfh&�*[�>6�*���b<BL�8%��W����.d�i�OsRU�f	h�Py��ߟ��� ����O��ş��v�9xl%N2�B��ԭ��la^]T�	Zr~�0t̫�J��C�L�y��o��nv�L�V�쇔�:H�U'�:'�����XB�5��ϒLP�4t})�t�d��L�K�6A'~�ɜ#x6*�-��������dx 묂�D^�?A��DZ���MX���ch~=E-ҝAfG��R��K&�m��m��7���d�3t��|�˶�6�����
u���P��cT������y������x�ۺ_�e�G���6��* ����-zƽN�k��[�K�O�I���4i�ƒ�3�����OG톻<�G�U���Q;�����f����;} A�[>�־��K�d|(�$����	�����op��X%��m�v(��j2^�>9�L��A����Ak��7�����_w�6���jܿ���mL����*���㆏���U��Sz�.� ӓ�02�K*7y����&�70���Î+����=C�/N�k�<B�^Ĩ��r�p��ڃ�8<�q-$�]K7��_3������B��-��<KBGzwpH��? ~�{F/��#~>�yw�`/�5�	T'I{�K������[c�����h�ؗ�2�RMڻ�D���_>AӡCQR� �v[.�`RV2��7�>R,�����V�~Y���|-�M~� *���I�x��D�$DS��P�dé�Q�X}T4��9�e�؛�:�߳'����.��˘H �QE�Z�L�Ntao��[J��<o@�R����v猞Q��ek�THo*���{�3:�<�)�ؒj@�zm���lP�8�x��	����@�MlL��bď�O�|�cs@�����4C����'���)�Z�H�Z�&1=YSY�q�ɻ*1�N�sf��d�}�9�21<�FEU�]�˕�I��`�t���KƉяԘg��m�ZaQ��v��e���?St�78xF���Y6)Z�}���48���أf,��eTq��Z���<,�`�D���̐�?�}J�
?!��y��)�;.�O���t�^	�`�܍yr'.	{<Ɯ�7Ahg����=H�o�5����8碣Mv��1�C�
C��໽ͽ�����h"-v%4����s�	�1�	���k@�`�.��)��"x�O�����������
Q���ܢ#�u�e�^� �J�8U�� �����c��ȭj80+i2�V=�M\׆J|֯��:���M�@��$�_��s$���2�h��q�;�+�eH����������E�	`.�-'��<�HU��^x����T�s��� u�/쌛�U%�rĞ���{z&��,�ቜ1����	�Է}�$Ny�%���++�!%�t���.rvcy� n�fK��&i��h���xdR�,�H؃L#�FbW����t�t_tg;��
��#Ĥ��-�x��hg���FW��i��HG�G�C���A�N�ks��祵5�1����ڻ���2�_N
m!lې�����OV\��ݬ&��y�5��˼U����c�n&�Æ4�r�6�h��9.���܄з����+�J%ny�� ����|�
ֿ��B����o� yz�Qu6y�	�&EX��ZKv�{��{�i$YְP� ��&ZB�Aݿ�~C}$�޼�C+�OD���%�C��T**�P��˺��H8�羬�-^G'�IǠV.X���3��lD�P��?��0�¨��@�������y<�@��q��H�v��p/,aü֨Vc��(Ft5jn� ��x������~����y�-�C��w��uy��O�L?vT��'3_O�aizd���C_j�=�d�\��u�s0���e�~1o�VY1��j���D�:��z����FNs =�x+WQN�C��`v䈊dpU�0ìwл��)s.|R���'�>�o�ZN;���Ÿr(>���d[���7&U������v�,u�3���N�"D�"�^#�G��qC��a�V�9�w��ȃ��Oy}�U$���:�D��>��ޕ,m0�!��nTׄ���F�w��ҟx|��5Kvѵ�Ɔ���xG��z�i��v�|�b`�(�3��R�ej�
O�Ϟf��d��N���:l�e+��� �
�"�%��'S8�WdȒ84r��Ƹ�ߙ�>�j��Q�~)0,��:���bz���?!�h�zQ1����%z2�~��2����t��9t��r��z�LQ�mD��7i-���q�ORT̀Z�Z�Y�8���S#���B�+p���bw�n�Ӊ"�Tl�"��AK��{T�mc^
�������ikݗ��)SW���Ҩ�u��6�w�0������6�ھ���f�(v��#Ŕ^c5�P�^��V��~!�R����V2�O;��c���Jϳ
G��e��J��M:[�t��O�7��{8���C�:|/C'��i��]�򄅿S��}i����Fe���IVΉ���K�ZY���ޑmsFT��U_�9M����Rz1#Yl��2H� �
I�D��j5r���K�LB#�
R��y��7���T���N��kd��D_�u�9�7[��}�p}�RP3È!��݄9��,X�ꤑ��x�N��ȾCٞ�r��×!ʤ�L�xn�[aUϞ�q�@��<\"	��eS�z#i}Q�'�z�-��v��ӓ��;?p���TS���I���e��oh��z5}��g�{4��Nk�PX⒮�1� u)k�X�0�4��} ���sE�t)����5�u�a��+����GO�,/:��H���*&@%e���"�%����Ǿ���].{9���٨��:ż����9�pmv�a�NtK��Me� �z��}�:�>��'���ƃ�c�f@L��Nv�_H��Ri\H�>�J�X��NTh}�o��*3"��Y���5�S0�g���So[�(�m�G�+d2!`v�^iL�2��"�(60�Gj$��=1��Ȩ�⢧��zۧ���;Ƕ�.�1�&��t���U��OrN{.S�	ݦ�����E�>�������)�>�b�~����G�<�T�7�k5{򨐈��5�/��K�� �>JX$O���,�Y�i�<}�Ѵk�~�yE��f��3�������2c�u�!�-�:��߽��O\��y��~���~�"��Ё�Ȅ$�R-Z���RF���[�2��,��(Q����:D��q�����L~=W�Ǌ��I��?D�ŨC���o�2�ӭ�[�F��b��Q�c�f���]�����k����U[�����@6禚�0�(�˒��@��A6�9"r�_d��R��%���v)�..�"�@� ���������L���ԷZ�;ک�C�M��l��/2PH�$"d@��^�� �?�������#��/_��k�{��t�̵2�t�L��:?���#S�W��yVj$9o��d;@��&��^+"���ZK���KX B�K�#���ʹ��C�t��c�Wm�㌚��J��'��v�`��O��{%��x0a__����`p�Ys�.��r�;&ʤ�~��@�n���O�*a%��еU�c�@'nW�?������ݮ�T�)�HR@�Y���w�'
�`q3�C�8�l�=URD��R�d�bvuqM18պ{T������T���:�6
�P5�d6�ZeހUwI��
4޹����6qK\��ùvP1|�
�^�x�s.�1/ʼ�ږ�!`,�<�J�o�<<��ƕ�j[��1�![�����r8���r6�i#R��g!a����3��Q�Eߙ�B-L���F���:r�%�I�D�����J�W����~����ɶ�B�K[I(�\{�ts���rV�M�HQ[��p��_�N�B�ɺ��Kd\�1�I��~Pp�yJy����쒹m�_�D�1�o�RA~�j�Z�6����h�fٟr�dy��j��=�>g��"��<'��Nxm�+�ځr[#��d��yhj,��c�&eUi�7������]���ܟ�����g�(��<f���ç��}z6�$�Ģ �| ����F�|O��* X�쵭H�%�{f����y(ő�����I0Y� �7<��9.H@�2�w��H�fN��X�0ug��c%�|�!C,�<h�Ņ��	�E��#Փ�M`n}m�o](�{�u+�َ]�q���G�<m�y�_:yUj���b|~�o3KŀF@�Tq)�$���f�?m�O�7�3)tg#h3t��2�Wm��<i޾�K�
=����;�݅q��م�B�� _�r�˯�����?|>��j�-�f��s��8���*�⶘�I�S`!>%�1�-��0>�#L_�dF ��Or]��<�@�,���G-��Dj��X���aJqCk&��k�;騪zi=���D �]�>*�|DӅ6΅Ǧ}Y�.�o�V/�� y�Գ����������H�Jt��ɠ���9���#���m�sӉ-��]D^dի��U$��H������_����k��X�ej�͉L/��E����h<m��/�!P��z��k�JX$����4��Xs���4T�A`�J1U!����R��F|G��A
1MP�797�ϊRh@o罢��fZ[���)������ �Y���|B
!Y�	%nk�H`.�`��\�h��X�!ҫ���Y}�{kܘ+*aI$���Uf]�Q�F��>��zEWT�������
��	��0I�h�^�cň�c�3ag�`P���2BV��G~�{��L*�����61r���.����5�r��b�2��O�:�����J��N�?8/e.�;}U�p� �������|��B�z��2eb�Z����Ȏ��T*�}F�-e�G�U��,��в��g��i��^� ��S:b����}L7$8���S|���ᓚJ��e��ч$��"ui{�+q���q���h���,5P]W�d��Χǃk����Xr3H�V�yv�a�<��g���5C�]R��K�>ً���|ti}C��7��$B�h��iR�Ȁ��va���/-��'�7GkN���j�C���q��ӣ�R�~Ю�1Ź4�[��p2�c ��J�ɂ�?֐�|r�����Uc
��k������; N� �L��5�����]��۞���a�z9w>�]� ��ߺ��&Gj�k�F$ѝ0��d/eB�O���Y�,/�%���ݵ������}�`vLfT�P��D�[�TA7������67�U��)�����i.3d�a�Y{_�r��s;�ڈ�K�Z���UH��������T�=5�Nhp����wXlxVHYEB    fa00    13c0؞3�~�=Ƥ?��'�\�
�8�!���Q�R��E���K������	z�u�\��|�&S��V�ߎ&�a�������ꖪo��on�/.�ĿFu�h��f����>ݡA��&�K�(�����9�	�@j[��bV�)�y4��tY8SĮC�y2>o\j�ىs/�6��8m��R�6qO��4sV>�Q�U�e�CUb�u@�����=^d4޸OD��R2��[++Q�NR�Wڤ�Go,�g':��)��	$-,e��v{�Ґe��/�.574�
�oX_�E]����	m	��G`uG{�잘�I�H$ �f�e,@I��^��	��k�F����Lݫ���u�{�
 ��������Sf���â���g3\�Ey�i�M�]i.J�(T�u
��t��I�Dߵ�m�"�I��h�m+�v6��Z�[����Ӕ���]�a"_T��Ynge�A��ѷz>G�؆F�����:��m��� �<ޕ�lsc���W�B�q9�E[��8c�-G�zͨ<9���g�ZbK+Ѡ=.RE�����bs=%�"�=z,d��j������c�ʝ�@�+�%��OI	��j�Ki�m����;��߹5�����V�SҜ��6)�4r �xȤ̮`�B9�_I!n>m�g<aՋv�t��Ɗ�C���6pl����h�cs���%��W��&���=t9��9Y5�M�~=ܹ���(�FH3Gq�E\�u�82�$,`���]��e�Ԏ���9}{�:�ן�&��u~�M!a��q��)"�*Qb���������ҪqǢ�e崣��d���2�4�E����`���܀�)�xH-�cn�i�[56&ր7��o�ժ{�3�n�s��_�6h�\єbp������E��6W�φXI���S<�l_\�%��Z꾌�D&�`������"�A��]��NR�y$V�q����`�\�[E�4O��Ʒ�ps�un�2O�[�t�	� 4�͈����wQ��؆���<�VS�C5�� {jIk�F��0BXQ@f:��99�q��)���D�NY,-d���v	'�P�j�g׆� �f?��N�\nft ���-�U�Lf��hB��N�rd��[B��GM��ݕ 	q�/�bė'�2nMC��L���4�0�v$��IF`!w��:�Έ����t��)��v虾��#���(���t+:V!��gs���ע�*�AAf�.E$HL�r�h�H�98�;ZS�kRѐ�>$U�}v�@#�a�g��� J��DoFy�-�[X�ʛ*կ��7��g��鹇�	�3Q�x���Ѳ��o!�5��t
%�T>M��#a���C%x�ԣ�n��D�������+��ݑs���ÁI-�V�����������A+].9�+��_rMv��<��kCm�|S���A�B��#4Y�����5�#�L���=�GB�H&&$�ꞇ9;X����xgi��7�%��d�2� m��Vb��i�|ɟ��z�w�ȇ��������9���O谪"h@J�(7C>+0<�ʦ�j��Y9ًƨ�x'q�K�O�Onf�vh�.v��Q��U٘n�3V�
�FS��!#��t��'u@@�vg� 6	+p�|��ծ�N��w�Yd��&~�p}�&�� jj ����w��9����*8����jJz�+\M
�8�&Z���d�<Uȇ����O�N8�Lz�̉Y��?�6��~o���3NeP�B�I���
�x�!ء����gx�;v#K��G��*g�n9��+ԭW9|�v
�B�J�7-��p�^͸�Z���-p�^�/�Vg4lZQ�ދ�R��㸰�7jH���h����RA'�A��<��<��]_���������5�9�v�a�`�W8h�� ��2�6�L/}�aҾ���"ă*�ZN�o�M9�������`暄�������F���IYoi�'$1�]��;2�t��������@�_h �d��a�Êm_LU	��n�d�A�8�-�Ff�8��HK�{"J#\lԙ��Ϛ��P4ރ8�H�\U%7.�����=�[QV�OV�#$�e�M�G"(��M�;G;%�"��.�,)&��c'���w{�Ɵ��>�X��*�5��c��Z��i&{��<^�������
��%8��r�JX,�gzm���}�+!��E2;]���9�g��&�<��x+�%�]V��K��ȎKIc�A��Iv���3�fZ���b-0Wx�8-�̇E���4�uW./SL�+�0��������w�!|a�u��?��cu<B���SE=��fCm�����:���
U�� ���.lei>jq�{��(�1�
���=q��c����ʦ��ʉ\������|J�9r)i����9�}݆<��W7=N�� 4���n����!g�S�R��9w	�Y��ÁH���<f�?_>�M�����+�2%2L'ٰ����!f��d��u/0YPL(�gv�P��,cb�U,8�s��vo�����"$�jTi���F�[8���idIT�1��H�wcz�.7jr`�>o���# (�J��(���HAV9�����i�,�z�6�Q%-.�M�MI��n�`����n�%�IL�r݅��1;��ׅ_�U�������l1݁�����\������} "�%��/,ͼ���7]u�_�`0��S�Y�#�����߯�_m��iM�~�E�t¹��Rk��"�N/��Y�W
PF%�߈y���K��P����.�,�23����C�j�G��u]�S.����
��=��Ld�td��Y??pϭZж�pRd^�p]� Rʐ��{�ώ/��<dm��!A�VI�������
���t�߆���!ĺ#�x� ݫ����|�8{��O޲�����O,�f<N^���y�������`빠��W�
�ʈ���Tr�����m��m13�<lUKK�L6��`�$m�7]�L�fN�O�A����s�p�������`��F`8z-m�<�e�<�o���,}�Eމ����뱣7�E����`�9ZZt��u�����X[V��>�y��D��q�q�a]z�ѨZ�d�/�s@��-���pp\�]<!�DO#+�'&��������<N{�i�Y�O���ax�һ;�$��Ѧ½Iͺ5�7p������w�~>-�wf�2vPtFO�c��wq��w�NR�mb��
R#U ��qI��P��G�}�9&	�O��ױ ����%{j��c�G�y��l� #OVM���q�ֆ3[�5�x��YF�!�{3�N?�<s��J|�jt#����i��Ha9��⦭�W4>Z���'梹����Pyb����ot������)�ޜ�#��I��-^�fb�#d+�&����c0�O_�ݘUsD���?A�[�ڠƍuh�����U�p�����e���f�Oԡ*<�iL���D2w�R4}H8�-�+��V���\ٻp��Ǧ�D2ssK�U��`ߤý�<#�zd��l�G^cl�����qE�(Y��/'�!�.���C�|�4,�kU_��Z8���[�`X��X4�p��m�_�j��'qG����.�y#���K�[ĎE�x`����DQۄ�? �g�L	��CT�ߏ(�H�,�$�Ϝf�=�6Y٧���zj���Y�majv����a�9��P����X��k���uO�\?4:�&��߇n���I<�p��y?,�Uub����5�Rm�N�=
�?�%3;f0�P�y�y0�isG���PL�&��k������7/{�kw۷�Z;�I6�|����{"#�tbw7Ne�S�	����q��_8��}��X�ۤ��������m�M�@X�O$]o��B���,�G&�ٕ��H������.#��i�W�D[�w�}���5=.���?����9�b20�m5 ��Ĥ�UڿX�k�4�b)��|YJ3/ѯMG��R�:x����J�'��M%���]����V�k��W	�O��$��"�&y	׾���,��B(y�y6\�������^��J�/�7����q����� �܆��A�Svi$�'�8�����!,g���D�5z�.F��}�B��RV��M��/�Rꚵ��^����s�WLGb	��%�󖅩����?��9�<�T	��7�9m�f�����y�$�1�Q+����=�d�j�S&G���b≦&����V�8�{t7�#�'*�3h��[c|Ma��_G����@��I=��+�b�ud���,	������)�;�p.i ?��Y�VO��f`��Lk듚�'+�\r�����������>6Q���pEՙ��w�6��Ml2����H�/�P^�W?;�ɌT��	�~dr�=H�jɗ\��7���Ɏ-���  �h߳cQ�\-�t�|.>)g��̥U�`N�ɌD��)i��A:&5pc��[g��NZ�P�G�{������2�� ��4�;7L=_[n�o�ג�������t��A��U�g�$ر���r7�bz��i0��(�]?hd`�Mj�í�.�>I��F�3�k�ڗ�����C&�?���bF�v(��-����`�p��Ȅ�Xh�܍>�h@C<�A�V3~: p+���t���P������m�}�-׵FX�z�SA��c aU���7��9�y�1C�{�F���H�ī��xnw}�M%J	mu�"׉�8��TN{�ɯ�]�����sJL(&�A�]����sT��\ų�`�L+�2�?��o�FjĤ[��]����ei�6D�	66Ѕ���0_��6���#�E *��&��]k
a�SHe����Z �p�����Tr(���V�|}~>p6y��0h�����)����Q�V��m�o�V-��wCn<L�x!o�@m�..�@�=�ik]/��'�W�uDU�54�j|9�ԇ��Nڻ�$�a����2�*4w7�l����c�xǓ����$��s��u��[*�׾�K;XlxVHYEB    fa00    1750���Q� �M�M=�	�u��`Vo��k/��H
�C^�$�M���ҐZ�7p�t�����A�U��5@����T���f�c����c�>%���ڴ�Yn6�B��4Bق�6�E����0��A�l���_�T�g��O��C�٪��*�*��Z�66����.�..� Ҿ�y"��ߞ<��3Շ��_�$qZŴV�ژ]����Z�PE���U��V�&���E்$�_ZE��u��W`(��F��ٰ[<�[�p�N"��3����Soz��B��B�-��j	�H� 	�t�N	V�g�tG�k�Z T��er�Cܗ��"��M���1���~;���j���&��<��qdJ�ü�>�#^�#�d�fؗr�����Ǝݲ����S�Wa[��w�Ia����g�����>k�t	�2qlil���*͇�tƙ��3X��0���|��eb�hn��:�35Fܹc���Ѷ'����o<F��ԧ�f�EK�d��� ��!n��m����dN#�H��P���ATf-.�.�3�0B��-�  �{����j`�³nU�~7L��]�n�x�ق�U�iA��
�f�j�SP�Sa����4��ɦזU�w�nbp�\�aX�3�2�kZg+?�`���
�s��}��Trg�����z�k�Ii'����K�k�/�T�>I@f�$��˝=�[�cb[=��Q�#�C�Ƃ��יI�a����[s��D��2/*�eQp�Q�MB��1	�"Za}���OqdB������թc�1�9ڣw[��|�ހ�
_j	�G��3m�(����T��^rc�A�f�*�*�����	$r�F��h�0��̷��֍�#�]�q(g�$�����n�dsPCc��s�����W� ��tI��{��4<fښ���*����8�C��x�q�ö�@��A[Ợ�b,��³�l+��7ճ��mx��M �5`�P�&X�T]���|ȹ�RoE�2Ć��h��r��3�'/��݀�S{솽$���Z,��~dƭR������j�����<¿>�o�99D�B�X$���91���a	��J�����Z�����f��Ŵ�^�a�R�~�Q�G`	X|DZcM�Й
�[�ov�}�W�>�n����E���!���.E�"�/J� ��L�����Y��r���еh�Z)߃
�1%B&�\W��Ys
���x�/���d�5U���8����a��x�*�K�9#�k@
� ���J,0����S��� �ʄ��k�h
M9�XvSn=0k�C����U����J��5�lIC4z���I���>sT�])����jW�\x�F�"w0N�s�B���Ap���J��6j�_">Z {D:��Z|g���0��h%��,ˆ�>�
�,W�ʶam�)��^���T��n���j��.˺�J�xos����D�M&TD�ܧ&-Mq��Jomun=wA�.>?�?�B��N?����_�/� �b���pV��"H� �O��\�i�rj�F�=6&���ɋv�R���kK����Kzp4:۔jΰ�v��=���p��
�ң6���e��ne4(�����H�X0%�E����26��⮻�KW)p AWÌ���A����N���6 I�۟IT�1����vD�(�F�J@�ŀ@� n� ����"���~�O��5H��27f-���-���R-��%p>�amp���������r���8���CX�U��v)����F<����otL��}}��4=��2'R�o5�؝�Î�"riU
y�R��h~��D����c)�	@�Q�~jC�Ob���^��:C?�ը�D1�ǦĂ$�=��N�m�-@樂Zd�7[�3^W���_�A�q���$	,��#H�J��tt�W��!���(��a�cΝ��r�D�����Z��R�9.phӯ0��ت�	4�Or����Q���-��������e(��7�Ĥ���G����(�< ,��~�F�`D��W�1����#�=�>�R%r��t ������Ü����u���?h�w�������"B4��º�ży%���۪�������~����[q��9�f� ��P��Y6��	Z��Qˮe�H��Y۪�mM�dCT��i"
!��?c�\�z�_�
��{	�W2$��5˔��KZbb=���<*C�t�Bߘ��<w�
�	FY4d���$��Q���Iƻ� �q��R��K8j�=��A�X�~Қ�1��|x��������0C�}�#�G�8��[S��#zl&��?�zlmr��f��'Xۑ�s$�D毳�Ǩ	�|��e��s��@����~O��x�D�Ѣ��f�?��B9�̎���rn��B
0��v�`�߃(k���F'�OW�"�R�3�����/[� �il� �)���ɉ���L�c�XC��x��A��,Ȗ�{Z�*���s��z�J!p=�D-�������8c�o��� �K0n�
�f���cg�0�d�?���BbWt�;
5��53~�#E�� ћ�HqF5B���`���_v�T5�����\W'|���\	ދ~Bd����]�XǑ/��\��0�k?��p�@3�A�~ɝ�±����w���}� �`t���ܷ9u�tS�@$E�%?�&Jdr�.*�_ct����X��Y�$���͌] J��Q��۾�@0PZ�B����4�V���Eo���,Mi�KWv�^�E�7�@������F�'mO"W���_p��(�"���/�l��"D������ub��*�_1uX�����핊P��KWH;�?�ʞn��bR�8/�4�퇣>Sނ�E����g ���&�Z��u�x�ֶ���$ħ�q%�T򬊁��X�b2��Ҿ�w�c����;����Z�b�5c�{]$�b�ezEp$�L�S�-�W��PSNCR;�Q	�.�<-w6v��6M��R�Y��|��<_��U��^%���"W�6�l�Ǘ��pS�.��TVZ�ܳ�
��u{ǀ�������������BE8��D1)���҄�YS��,W�t��.�H�۶B�q�����Oz�	��X�VX<�8�Q�__��5��	��[r�;�p,�q�s��e)��V�(-�EÎ�X�>[W�����w�X<�D.�.���[��nV3���{���ޚl��s��e�9���
��v������2�-��Pg�Vv��b�	�S������b�?���Ӻ�t�uS�Bh� +1�81�İ��1WJgB.���M���&'�\��L�]Y�O���z[߳h����W��R�V^� b鐡���ց�b˞~y9B�o L!��X�,��3�0�/VV�:
���m��|! ��Fj��30]�&����X��g�fo�Oh��7���� [��\�Q��o�v�A��L�!�����c���s�Ge_�S�O���z�i� R1�;��<��?nz��A �����������a�k�*o'D����ٺ�$}gN�R	>w��݁o�%HL�>�׉��K�y�$�M�t�ͼk��u�aj\^�Pd_�(�
C��u2p�i�[.�E���;�L��bx�����!"M9�NGյA���W��ޫeSNͧ�$
����OYy�n�� O#�Y�(�Ĥ|{�_�"\"<��2�@���DJ�{J����?3����Oa�w	[&���:��a?ʎ8��nM�l�!�U<u0B�l+Dp�ve��|=^Z����ǟ��很���pM��Nn��-+f��ԩ�6ƕ�����v� *A\T�ig`�-����Z	T!7�!�BĤ<�:��a���.y���zi��F*���$JEk#������C��-��
B9͢��R�T�o��~X��ʭyM]��T��[� d�-^�H$�&�3��)B[��ە������=EӦ艐i���A��S.k��A�>�Y��o�\7��gQf|�#��o9�JUf�J��O�fr)��U��W�9ěLG�Dtnvm��>AZѼuo#\��?=F�>}qP������"t��NpBq!��^�Բ�b���lQ'��!����T�:,h�9�l3sF1�+�� ��$א*�o���7��JJ�i��iA4�ƿ9��QVa�L��v��L��)�߃����~E�t�
HUʬ�ء$R��~���t���^�<{w`��H��}�����P�����Hm�7�Κ�:*>�I,bc�
�v�G�z����/ �pX/??<v%�����C}��`t�ǧ��ŵ5�9$Q���Bj��x��A����Y�h:��7�>����v�?�56��~Ĵ�Is���:@���2 MqϠ���_#�<]���
��J\���Cth�f^����~�~�	_�b p_��4({EmE��$���|����;�#�M?)��U�P��:r�>	y�4���gԣ�;�*6��� ����:���\���rߕ)׈ɲ�R��>+�ܼW����#��p����D}N�Q��6V���8I3��$�&P@θ�6K�T�nj���<�=���R�fe��ן�S?�|�5��>�$��d	'�_|�c�U� T&���j�,�}��ڹ�R����>2	svB����d�TsK�f��q��dc�1�32��:V�����y������s*�"-gW�C�6� *�e�-x��k�{�X򾬱	�Ǽ�W1�����v�&ׇ��B��ً�+<{k��M�Q��m�ê���z��Bx6� ��ٻLbve���YIM~!J��38jͯ�.y{P~�P���]]���b/��� �i�������.ĳH����|x�wI¾�<ϙ����D��T�j�?P��j�e"��*�<�'�v6˭m{`>���fMՄ��F�FE��]ޛ�<[y�D:3w4Na��Bk���R�i�U��w)��8�U3�;|M�'ǒ�M�\�1,d�N�j���7���qU�����p�y��g}G�7��>#���鳢�k@G4ג-܉�Ӌ�)�)J@'�!��{$���9}jV;jҪn��
��Q��a�&}��������8�T�	Ǣ�s�bt���#�k��5��9�ɛs��``�Tg0�K&lYs�{�oI`�ѩ��;�e$���M�W�o.��h�6!7a�L[�dM�(XfbsI���t��+r���v�D?g%�x��+���SBT���<���� �䴴��T"�W�����E/��ɨ8栄�'�%�_��%�1�MxJ[�HqDD�Z�DN�Թ�h��1�Ew΂FIL� �0U�]@���w�O�Q��[�Df609q�1ҙd�,����E�H�Y��;��N��%���)'��r�����qe�$r}����&�Ad�9����ñ��^�4��e|��;��o��qo�����|rN�q����sw��Tk���W�
g��X.1n�7gmN�a\��)��c���F�kȞ��HS�'��C��)�����f��&�Kv�xyZ�y��/�nmʹ��hǋ��G�
�ne�"�\s��X<"�3���!�H�jj�g�l2��
�aD����Q�Uh s�U� n��N�3Ux���n� ?���O����fr�Mq������c�L�G@���l���u+T�����uB/Y����0���2���@=Շ����kʉZJ}�@̑�~QE'�A�Z�ST�k�߄y��Ѻl�H���6����l-K���K�1��p�]i�Z�A�3U�0a$���]I9s�mW`����txAro�Q_�?qP1'<��+��?���DRt���uoS�m��(�b*X$Y�+�����话ݷg��XlxVHYEB    fa00    1870�q���tL��ѵ���I�>��̅���}#]��8�{�&�����߭w����P�h"�z��8pN�ߨ�r�}�pX�NTy��g ��#'�ſ��H�*r��z��b�v���k�,�✤�F*�Q��xm�q�!��%[�FuQ
�=n}J�1_k��/�Xh6�=�(���C���5$�$%g�k���DI��X�9�ҳ8 �M2T|��,���V��h����%2��R��a3�$vͽ�-�>>��=8�����i���c�ޗ�r�1P:�ʿ�v�.���i�-6��˿JrH̋���ol�(�7����~":�z$��i��2k~7�
����ۥ��`���w((N����ډ�X2qq$֏g$�a�]n�� �T��CM��f�8ϕ$���Q��iY�F��E߬�o[����T1I��J����莧?_u��<l���{d�0Sn�8�Ng���(�MU�����ډuF�a�
нv@�����7�m�0{}Cj�p��>����,�}1��ek9W�-�X#f�M*]�s�(G��ܴ�����7, -�@��
t��X�zMc��w9^
z�D���@�����+��N'�sQ���U۷}4�B��%)ݰ;�`�'�,��X���I���AQ���x�k � <W8T���K�
��n�#5�!�z }��U��CP�sw��O�.�[�]i��v�`=�(��l���pm���}ֶX6�Eru��Gcܾ�Cz��PZ��[�$�э��q��j�Y��2P�Ӭ�4��
� ~}�� �Uw@Ṧ�h�U�y!q�� C,�6���-�)�E~!b�w��l�̗�^�*������^UP߶CE�Gbc
st�R3)&4水w\�7 :�W-�:�n�Fy�Ao���lb����3�d�����~;��`�:���V���� ^J��U8�E7�k�͝������'�����S���e����e�
9����ŉL��_������X�(���N ��_��9��k������_$bj����K�Ċ��㓯Ar�J�X��Xh/M�T �ݲ=�I��p�R.a��tR��,�d�m�R�:<��������mA�/p��Z�T�I�]g�l��MՈ�K� e��������b���a�j)
��A�D�x	ЇV��<��"�-u�4ŗ,�8�0�Rvv9��[�zTw�dR@�ë�f&ѧ��/1D Nz�N���Rt\���퍭2���0�����WBI��uU��Q��Y
�uR6�Ð����o������t���Fǻh����{����(�~?�U��Ϳ#��o��<Rl���-��I����@8Y��.�d�1,��u[��yE�7wKz�F��d�r�Hr�\�S�#I��i`��9���߭H૽�,��an����n��q�B�� U�!muV��T�����������й+1�93�i��� H
�^V&�0����I�n`=:|Ԗ-���!XdT�sul�I�x'�X�-�Y�nvV�"dU�00υ"��3^���k0T��H� 	�{�������
��+X�]� �=��Ǟ�q��y�>��ܬ�8
̈��u���O�#��*Mbj���� {�ܛ��Wc�?���1�0O&k8�_��T�6QU�'��A�rQ��A$ƚV:���y�.� !�E��YE��$#�R����=��@�G<��?��B��L����޳�/�W�rd(>�\0�_�d�v�_�e�щ#m�\�:�i�H�7��`�	���?�������?n���2�r����m��~��^�R��(l]Aދ�.+v*H������qc��7�KT+� ~*\	4�d��I����a#D�$�����:y3~�3�OQz���Mp�~j���+V�t�`��0�w6��]���kҩ�'~k�D��K����(I�}L4��I��e����D�1َ)Ӄ ���'~_5��^����,	D����z_�RB���P����i��4���K��	c),rm��B?0�J�ݩ�S$֮��Q7�X$[�t�i���?u�\h�Otؒ��,ݏ�A�[e�Y�l��6�^4�����t�F���n��1>q������Q��3/�c
��q���E���'�{bS�n��<�$=���_��եCyEc�Yvn�<��Q�����uRp�W)�a_�c4d��0w��8NrcW:ExB[Ϲ�T�D3�k;��+Q�ղ�?&^��i��]K���������w����FZ;0`?�!�R*F����
�.:7�'�h7�\s�d�鮳Pn+�e�m�6h�u��L�us�H~�&gE.�D��zdnEH^b�	��a'덱�_U�M�a��4݊sm1[�p�t<�/
A���"��|�,�T���d�tN��Q�3���#F�#?�t���d	q��YWi�hv����`�0(o���/�>�QiN6������r�dM}OA	!����g�)r����%��OS�Ԯ�X���mG�\S����h�5�뱕�|��L��
��yzRw�)�W,��O�M��h�p�N��>��L�]i���f�Bl�������G�m��eG��0���~\/蓙i�N� Q*��	��4�ڨd'�w*�6F�?2ZSi�.�;d,<7�g�D7ղ�&�?`�S��5�mi���ji�ְIW6��ێ;��os��J"�廍P
�
y�Ҏ������_|��_��;c�m5'���� ��J�?{YeLH�n�n$o��H�� ��X[��n�@�&I��dT}Tsg�/!���S�1�$f���P���,��	�Y5R����� ;1o� �%!������T�mA�.���AR��9<$��r��Q�u��fa}Y	�Ln�r�Sh�M�J�jLwQ�6���Z��z�4�̥纝-���Z[�z����LiΞ�2��Ypҽ����yJ�eЊX=�Fފ:*L�o��������],�礆^�.u���w,˪��ֲ����*�j�Q,��:�'�4���`��}Ư����1.�A��>�Cf�	���+ӝ�S��+G��F�V�W�Ǌ�eו��'BR�XD�>��'|�P$Z�y�{�.��\���T��C@�r�N�����9��`�=)q�ĤQnD��Q��c�M��� S��<���j�g����Íp�d(���/S�{�l��,��l�
>ψ�%�UБ>�;�s
g�o���R[D��E=p��jE��;sԄ��n��h��n�:��h��	��˃r��
s(�7�R�}62���z�5�����Q�1%tm0�p'�����A��H�G��(Ӟ�W�å��5������������sst�|�����e���#�,��Y��X}J�)�+�}��W:��D6�#,�ص%AYM��<�2�1��vM��|�H�ߨ7�/��<ư���Pxጥ���-"�C}���H�����_�K/e)7��J�O�7��F�U��`����VXR�܀O�as�xLp(�u��V����i�0�Fw��Ǔ)?��âW�ּBL
�%�_�|����cA��ܙ״S&��X�΢�(�D(�!Q3�S��g���C��0�.��#�$H�1������8��q�ެNFD벉=t%����\��^�=M/_?ˉ|w�;�&
+A�����&̀��������>��O��-p1�RoE�O�4���7ة��^,I���kE ���H�"r�\�z��!?�prm6���/_Y�sE׬��k�ⱘZBP}��]����O�M*�R�簽b�Eq)�b���z���I��F4�^1}|�U>9I��>������G���#'_�9)<n�1f,QiX�R�P��b�0S��ۨ������y֖�-�������\rZ�4/�䇽��OKR*�Z��K��	��oĜ�
����ޣg�B���2�C^(8#h��YB����2$� ����9���|���:�� a^�f�y�w��3�������^i���8��l��w;��"�U��Y�M'MeJ^IQ�!(�RL�����̅�Є1F��Վ_�Rя���l����"�V�q��sM�։��)�|߫�\���aౢrS�ԁL��S�l�����)�+V��5�l�� %�Ǔ�Z:m��C�J��n�� Da6_�L�m�4>�@,/��0+B��Գ����D�(�����E�n.@l�V�"��`�h��H�]!}�UW���)�5w��_����2y�jPY�C`e\��;�ש.�����G�Λ$�wu��!]|N6O+���kf纹&>������d�`tw�)�Ay�fZ[셷*\OIET�)�J��ྶsQ��\m��T�+�Rj����5'�1�8��wd��Z�k���W)?�?�
�1�6|C�4e�ɠ[yi�_��-~� K?O-܂0�iJ���t8��35���e�T��}��;�Q	�0��V�N%ī�ec�$՚w���訮O�H�E®+=�>~3yI%��ɍ�p�hB�n����w��[//7��겦��)��x^B���@�d�xr<q)�����ŰwV�0�Dӟ Gb%R��p穂��^��ݗ�N���1�E�cF��� ~��1��G(%]S��{�h���ƛ0�����L��J�KWK�}멺q1L��<���ظ犊*\Ӎ��B��u��WD�����F���"��H���;�|�{�Û��q=�N,*��"�#~��>�x��1d�^�Vu��1NiYBe&��8���,��"@'�B�f�gM�����C��<Em*6�A�qy?R����P.�q,!���@��'�(W-C��V�`+��qN�!��hB�Rby�����.�7�{�x�Wʊ���.��[.�tI�����C5�p4�p�����f�pH�5�w��ӄ�08"5΄&���|π�zD9vc(���i.��k�fc�Tă�T']h��������|d���UH^�&�2+�0O�}W|`6���x�CAq(�̜����t��i�9�v�3�N��;�]ʴ�q����@���n� �pi�Sl!'�N����l�`^�(�Wy�Yܧ:��O'���՜~�{��T��?ݫ������-ș�:�'�7٬:)o�.Q��DSg���#6$#_�V0͓0���ލc�H�:�Ә��e�P�����$�g�F3u�W�J��8um`0�-�t��'9�T>帚H�uG�� n_�m��7:�����2�ہnB/���4 ��oЅ4�-Va���
C��L�tV�H�0"M�� G?6]G� XU	8z�FL���v���u� � �N�UMkdDZJ�k�6����HÀ�Uz����N��H9~<���{}���%3s%�q��=mh���͸16�������W�l�L/�w���,,�]�9"@���WQ
�W���#�.T4w�A����ғU�-��������QK�d��0_���ܶ��cr��T��6�+�Z3��bt�:N�]ԋ�-�����T{:�ۥ*P�4�N0P͂H�F�`Y^��.�o����NQ������a�=����W�cL���
�
^�n1u����Nǳ�j�݈Π��,�7�lse� �~Ϙ�!���b�&��B��%����z�G�[sDv5
Pvd�^$ ���\�(���Y-��@���';0�!I4�pޘ�م$�K�������g
0$T8cam���?�j^�&cTb�;���T�K�<�*p��+��X�g�\�-�+Ȩ��蓮iVxLlD�T�5����1gdwG�Fe7�-�{�{�Ri0V;�������ͬ��-��K���%ÓmX��>�j�EcR��Z��	9�h|�l3�Hy�!ް`�MNT���(jm �[�����]U���:�9�>U���|�ț���9.o���[<�e�+����WU�ļ��#s��E~tN$�д7{�����v:ɖ	ΣZ�D��U�>=�*���	+1�*��(����Ep�O�}c�i�2$#�\�,㙌)q�x���O� e&ip5�Yt��>\�l`��^�W�w�m ayA��-��kήQ���i�?$)c��#!dY�J*r�xͿĝ���M��PH��[������>�s����q�1�` .���Mk=�׶B�"���O��;�z���qR/�>2X�XlxVHYEB    fa00    1210qMt�4��CϾ����=	�� (���b�0Q��_Jg�j%��`���^oeߟ�F�b}��o�y�[A�谪�N6�;����> ]�M76YP����Yr��E�qa��0b�X���'$?A��~��r�!�����|Q�a�ZN�����.�n'@u_��N���|��Nd��F [U��=�qk�U�0�����wO޷��.䌇@6�()į��K�i�� ������TO�j[~,g��(��(��U��Fu��c埙WAU{%Z+�r^�|��o�a��`wW`:V�R�z,��0�0y�Uo8�(x��cj��yB���1c"'*����;:b	��ʊ�f�x���YQ*�_�-<��Z�Ns�T����TkFk��_�|�ؿ��7c�A���9HV7��Xf
p%����J��h���p�N�'��}��XBaR�@��mːZ�y��O@vi��;X��H5Э�Qߝ_Y��.<:]e��嫚�b�w�:�c���A$h��N����5e�lړ�J�G��s�e���U���(�mU�c�-���ϡCd��iH�ː�Y9!�+�
�ݩ���_5Pv7�Ab��Pu��M�&@ �Jt?������6�k{���9>CEŀ
�/+5�V���R�'�(��1{�&!�=���F��Ɣ�����&K5ᩔ���0�4/�&I�P$�,-À�Y�O	G����k��m�ȦQ��j�(�Վ�`wĥ�4�F����78��v{��U�ǔ�4h��w'�ܰG���/%�ŵ&u�hH�j?M'�7���Q�W��a��ñ�3���K���-I[��@`"9&�2��Ӟ:g��=ͪ)P�"�8דO�CY���L�����װK��9�fE��3���Є���{#�q�m�pn����H��e����8~ʶ��<x��}u�1z94�خ�d�3W�g��|��r�
�>A��m�j]S�BN�4v(�B�Ez8��þl�?��޼�q?��s�~�p@��G��0��o�g.~P��P	C͈+�J'=��U�N�+c�Bh-���J�(�g$�w��.sV��4�ȵ��e�d�T׌#�/��<�g���_@�5.����rB���ݎ��Ք�sg4Y�l�|�����l�ظԔqN,�HZ}vȒ�eҕ���y
���B�����n�'�?�~	Ӄ`�/R�z��F��\o+O��T'+�(��-l�y
�K����qu����5N��+��眉�ѱ�3k�����~'ґzK�nܬ���t����3�n%g�n?�ņ/)�0ڏ��c�>�E_��9�fCTݮ ��:�ۡ���m���"�0)��6!Ak(Y��d^�����{r�9�G�\i��)ѥ��%
@�M7]%��~�"?<�H��\�(���b�#������f�6)�!���+�ٕe���y���DA�����rb�M���iY�V�\�T.LY�"[r���&�>����0�#ƍ+2������_�l�v*�7�G�9Y�PBkܦ�q47�\�'��6�b���3�����mW�
iҰ��ʓ��#���� ?٤�Z��"�c^$�F^�ŕ�8l{�3Y����P�<gU{)�Rv#Y�bH������տ ��� �sI�L�� ýذ^uq@�����$Z]́��"�! �#j��b'i�䕗��$���Z �c��EY�j��9��`!�R%YsM-��\>��I�j��A�$�o���a�����$�LN��7�:r�m��G�x�"IF���r+�0�z�Z�+q��w[2Bg�u$g�ٸ?0��H�ű
�����{���~�v�pU��H��Ρ���aK����o�aU=��H�[D�Q���E
/�g$�` ����#���f&*ѕ�H�2��ILiJ��F
��Zq�do%�]��\������ʀ�X��P�dL�p��Gi���0)8��n ����X>�h��6�g؛@�X��6����ܑӀ�_�{"^c��\rz�VD�n�����
���6Sf�%��9�c���!*������P�g~0����ؒ��,�5* �EXe��~6G'�H�*�(�b�����n/��M>kn�V�z��45xy�-�0�~H<����QS	����@�a�B����$�J"(�iqͩ<�WGUoA,|��[�D����P��l�!G[��`�;Oڢ�]���m�/�	�DOMw�a1���v��P=���1xk9�����F�4me�St��`�z��@��ZT�RƝW~_�xX�	��Pwd}��m�����@E�+���î}�/WQ��~Ai1e�]��@�����&W�ŉ&�^�?�bY(Ыr�5��4+�P�7&h#T�/����Q=�?B�m��+��</�:,�A�g���I`��;��*E��u��5�-9,�U����U�R�H+w��]�¸S�F���j���G�V sג�?y
��ٵܗ���@s?���R�_��l�6u���zܺy��q�O|Q\�.x�%��R�"u�w��u+�S���[�*G$���kgs�b��k����=�j,(�y���Z]�AGx2�_��{���Se�UP��]�WxXF�L��E ����/��1��fI�ҳ?zD=0�<�~?��}o�B��N�=&9�ʤ� !m̅E�Z�cԗ����Y�ّm_Ia�����M��h�֧��M^�J_��G��٥��m��b�w�W���!�H�83ǻX�؟���n�e�h�"�����xÌ~ QGKN[�`��b���3���l��Ɛ�F��{q5r��Lӆ�\�o�2,[OIx�ү(�Ab��h�}�v�u��R�C�GYJ;@�U@���N&�b7���̨q��8nT�q������:�#$t"��,b;��A�n����
9��I� �?��#�=�s�񀌕�S[I�XR��&F�<�w�ͬ��a$K� BK>Rv�;�0� �nD�9���,�亊��{��*�U7���\���X�h���-kB�c"�����'w��r_CaD�5 ��n�QoT8�.8�f�<�N����IS��D&M�_]}x��
6^2���{`��Їb��^2�<�_�gj�� ���ɨ��J�}�P��R𣾀�$4R�=���9�B��@�S��/��g��R>�+�6�C)�o|f�%1P�&��� ��=���� �l�ѩZ��=�4�Ȱ���NU���r��X�{q����D%��$<��~� ��p"B+��H�lg�a��o[2��DP���a�&.{���p�����^�2����9DCp�8��Ҥ�&�߄gW$b:^��n�w��{d�ض�� �0]��Y�c�jK^�NXƓF�GA����k����s�e\�^l@��d�X���.��߮:��/���O����ɯ2F&�b5�p%���%�����D쪷w`�-��h

��! �����5'����*u�~(vU9WZ�����!��V�O��J�F]��kW����>*c�q�JH��~(���-��Kc�>[y�?T�S��2v��k�e�틎J�]�9�	D��y�nW)� ��q���IPoD�����$CRB���.�M�mb*�*�Q��f-�h�2|LƮ�3�a�G��U�ꭡ�TkK�m�5S��F��66�b��kՊ�i̗%����I��/�H�st�9l6�cG�[}����*���x�z�I�P�O��q�%�0v�h���·�c��ɋt���P� Y���5��N�_�((%�_Ϭm?
�[����5���6��� ���L�RS��o��)2y��a4{\���	�ʠ��}�@^�F>b�w��vݢ���l�Gdq�<!" \J45���(y|TL��}����CUy	�ٹ�9T�.�^�I��TϠ���j����=
mh��W�k��9d����rq��\`�������vƩ��)��cw��3�9h=�H-u�V?�8�$W��[�w��;)���Pʭ`ߍ���T,"W�~���w@'���~%d`�*��x�����P���fm�Y.aA0��R���6�Q:<\��?�ޥK���h���r�@��ɿ��y<��\pF�W����LBx��r�(���[;����2E����驉"����&��Κ&k���g'�6
Y�NIcr�/=	��pJX��\Dn!�M\�5�r�(Ԧ5�o���� j�4���],�A�����<$IH�
r�p�;<F���������dF�����h���Ґ���Av�@�V0n����76	���:<�ƅ�NZ	�3"?�X�( E&-�i�5����Քc֘����0B3_��:ؒí? \���X��N�.
!ZN�w[C�t����rm�4l"5�������_x���|�$�!��`�L�żs1��^C���M�۠���� 8<�1��˶�(D��D2������:��[ef�~�r�uu.�21�^���O(
K{���C���n�j�;:+F/��� n�ȭ�"�M;i��fj�ƃ������[�WG�覶ޖ�3tl����ǩ>M�59z�������	 �W�Z��e�ĝn�8r�����u�/Кҡ�40����!k�|$�=�&�ĠXlxVHYEB    85b9     830���V�vn|;�x����
U��#�.{�p�ۊ�[�>^�5C+��)�XFo�M�Bu�}�sF�a���z3��s/�K���qB;리�����^��>ۣ��t�cK��1� ૭Ck��E����2�&rIu�nn'h��].���2�	~ח3k�K��k��G��ynTF���s`-ڑD*4he��,'��8.,�)f݆~Н�G�g�Qd��y9�{ç��2 Sa�ÌX�t�SGV�����Dj�-��K!L�Z�&��&9Dh�܎��4��$�vW!/Ψ���p�z�F�O}�<䌞O��'o�(��=Q�R)1u����o9��%��r%��!��Y��?��ʽ�fo&���2>ާ/��r��*k���xi���o��2h�,4�ܠ�gP�W��\ZY.���e��T���,�í���@� A2�8-���=����R����g7R�[r���j���Os�P�ٵ4�,
ik���3�5_� y�r�2�>5�a��$�z�XƘ��vÊ�L�N�`?��fg��@(�J.�b�V�(��!\�n�#A��0<ثޠ� q�M�-C�T���� ������m�(�]���ȈN�����5�+ ����n��>�V����;�NQ �//�W�>".��T�1�U�X�#��0(���鼗Y�&<��t�#j�b!\�:'\��P�ƾFZv�E�"�z"�2*��BXZ�B��%^��ǆ<<��9ݏ��t��H�g��������/�$ZXӢQ/���/�$u�@�ﺫ�K%t��ʑ-nk�-$(�r�#�ftL\G3�
+W�g���!��"���(M���c���[*q�V��E\�H|�&`�mN�2uw5]^X�f4���.���j���M�����1��ͨ~�U��s��{r�~�U%5UM��©7�t�H���
�Ǫ5�� �����2��G4*�����(� }��Y�r7r���>�����3��o�����,C�?�3l����_�r0G��wr�sc����m�^�����6ݙqM�J�Ӟ�/�r�waAx�~�|�d�\x$�����x��.0Ve>�j�3|����3�������Sq�V���# ����D�9n�Z�����z�q��a��� �~��#���~�} �yC<����k�r���܊E��oR~��rG�*�b����Q�j2rAR������x��4џ0nh['ݯ�~�卷׼�A&���}����T�3����&�p�u�J>5(����<2Ġz0ؔ~�}ypf�q�=h<)4�������MXcD��7�"�k|��D��O��b�8׋r;[�e�oo#��m�Ցj��ͼ��{Z�=�F��K>cGVLs���ȱ&�q�:x�r��`azHZU[����v�3⧈���b��e���$��K��y�ش~��8cƨ�E�1����w�6);	�z�%LW���v��MX��3�qQS^g��(m��O}3i����υ>R�Uw_�G� I}��y�!^�Ku��G>��nr>�Nxה_���=�g�4+���:H���R;�W2À��L�>�ǴS�ɶAd���̚���f-Ɠ������.g���Ϥ���H��\��y��#���x�5#�nM&v}��So��)�ڲ��ѰA���{�޼�=94i�g�AG�Y3����<%�;�)�����������6?�́�~;�%#�<C���E��;��]fz|V�ɪ���g���cA��N���Ҩtܩ)��
'O����R����܅��$�`��Ҡ񦨈a����r$-�ɶ�6��S��e�2�߽Y\Ĕ���Ôﷅ�� Q�T�Am���q~l�7�𗽏��}Gi�%ە8KQ8v"y�
�*B��/�z���A	{�}��������^�pp��f״&B�e����a�$�P�hf�Y���z�����
3�D�s&�j�l�Њ�	��!{Z��B��
�=�<`҈}��'�DL38^���ҥ71�t�Ph���:Xk����6�\j	tPcH#b��mY>F`�L$$����