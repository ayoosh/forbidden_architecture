XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�z���+"(\<����}�����-�ڌ[�ce�N���]7�Q� ������-n �+�⪪�#A������;�أ���=�ჾ8�K��ed#@�M$��9g�U#=��������W<�r���O�S�h�b!F��@n��u�8oG>�����:�7]c��*0��	LD��	L�$;���H+�7��v�K
Є=�cZ���=,����W��+�.�͔�T?Er�"]ٰ��3�cuәGV�����!KF�
�=�Ȥ@����o�=������N^�n,�.�%XN�߆�� ��p��*�.�I��`�W�S�P�f��5����xv`��d�
�q���~E�=�Z� 5�|�kb������]&6��������T�UFo�gS�����gPuR���Joc��6��'�t	���͛��t�w>)���m~d=0~s��V�LeӋc<�O�8�����7A�����~l8�f1�r��-���t�⦽]F��E$�xIGb�ܙn��#1��3 ��t���bG#Y���U~��%��{<d�I�2E�����ȾYNkH�?���b�z;;Og�Ŝ��ny�IyP�5kN�C���~�!y)��k��y�m�H�i#�w�0N-E�lPTk<��%EZ͛tC��/�˾���,F����q�g2P��.��WJJ�6���	�B�fRj������}bY��Rz(�o1Ӏ^��C��E���Q(����ʪ
�'"S!2��b*�s��zyS�s�| s�XlxVHYEB    9de1    1670�+ï�b�y(���R"Y\��?�>3�f�>��UZ|�[���_e��#=���/(Ok���+ߥ�w�)��oh8J'H��!�DQY�Ci�ImH)�b�{��W'~PRuWE]���vQ3$;`�)'8�@��r_n�kG��s�@��eSY�l��O�����׀Twp/��4cel=(X� �U[U�C��z�"Y��"6^f�уN�>�b�]�섰��gr��H�{B�KO��'���t�x�|���F5��n��2�EzK�S����`�O*�ԙ��z�b��h`�3�K�Z�Y~T}*���a�YH,��@t�?���
�m!�ƢG5���M�"73�,#/��\�˔�D�8�Ĥim"��0��m)/����\���K���������!��%�<Z��r�� ��$p�5�"N}��#3мp��`���jf4���'6�=����x\!E��Zf���w<m�#�5aԎA`�~C.�Q����b�T�Vy��1shm�mw�P�%I���#�`�UyЦO�vZ�<�Y�z����6�mnCOeU�i��]��]���C2!n��wS#�	m�d���65U�-�tQ� ~H��D��拊��f���~'҃��$"V�����zRNA�4=D�E�Ѹ��ɹO�-�^��{���`�H%�cعk�K�)'v�iҢvA��.]�.z!,z[E�����e��F�ɕ��ӏ��6'�v��؁�S�\���@�4��U~o��|���u3�S#�G���ǼÅ��CL��=|�sm��%�t<{���?��a�6��nQj�g�3ƾ���nܯ�*�9n����iQ	�iDo��F8���JkiwJ�bؤ��8��
� ��0���k�
����1�(:�T�Ɂ�(��9X�p��Ѱ�%r�b����43w�}�7����`�}��	Ьq?2e�n��Ba�~�|��?�������g��0NU�������l�r�1ߍ���0t�)�]NcD�<^�.pF���F��UI 0
��=�x]nV��ڽEJ�)�h�_���>^�p@p�U)��"ƜB�-A$aJ��X_�:T���r�"x�f:��O6�bl0�t�_X8�x��t�#�H`G�no�&�YKMT�Ɏ�!�� ���P��KxN%\��E{�)��ܹ^K��Ga��p)�5EV8��>��VE˿`L|oEUu�œ�b�$D�'I�2+�alI�����"p���7��č�~~�4���.�*f6�!ի�� T3��W�����`E��G�-�.3��
�~ @CF���DT� Bͬ�Rd/$tU��Ӑ��`f�i�-	[/�����V�hS�*�ӄ� �)���G갿�����I�S�~�)�/7�=�w�
_(�_;�����(2�ϥų����T�㌔���i,ɲ��K�7*:Y�\����m_���+���#%��]7#�u�M�l�67�M�>t.������7da�D�Na`x�-�"yRʴ�����4���U���"�9�
G@b��-_4��D"[d&��k�Z`���ӥ���Űö_��.�R��l'w\sS�8����7���oyA|� M�:������������#Ă.��e��/GS�-��BI��޿� �;@�}�X������D»z�k��b��ذ���v�D��\6UC�˼ѣ��J(���_��������=���	����������n�h
L!a�f�x��(�m���SB��נ����%�~� a�C^j"������C�M���N�b^����1BJm��@:��dʝ�5P��g�}G�X|�����ԄUBAҹ���W�E���_�����e�����F���j���As���W��-����E�����7�� 6t���7���2��c��k�;w�L	��G�,;�/%L�b�����j Dp�����]�꾵����N��b	q��������R��m�P���fEV� T���þ @^��E�%I�ƌjqʌ�
���ݰ�� ����T�i��0{S��w٫҈}���߬�8*Y/)M�]6�I��e���R*2������Ο�2N���� Ճ_�e5�8u�HZ�� ��K
G�C���&�|�9ӝ,�ZeW�%�Ī�����ݠo���'YBeB�ɸE	��Q��� �����U3܉��Q9ԅ4�V_�������qn���zL���w0��&��	@C:H�$����۱&�X������W�+C|t�>E�?�8�.b�ppm4v����!}M �"h���?��_e��'*��ju�=u�5�ݳI�q#�Y ��Y)�ઊ���^s�$ϞrT�& )pZt�A5:I��FJO{�iX�� &	��yg��X_��q33���km�~�O�&����.`j���8U*�]�Ɠ��,�U�����zk��8�g�x��z�1�W��<����;��DTm[C�Wg��� /�z��f�������H|)�	k�~����K�o�()�[}�O�O`'s����X�-�*�~l��#{�^��G�H�cu�A�P6s]���2��'��H�{���!�$�?1a�<^3=�
��
Q�7>N�*wI-!�U1e�Φ�ㆈQ��7p�-��4�w.B[ւo�1[5�6�l��W�r@�W1�}Bo(����ވj�Ģ����R3�����5v��t�����a&�݊jz���"X�{So*kD$�kG�4ۨ�dSh0�t���^Ì,M\'�^i��A�����k�i9���ԋ�ʓ�Zs>nLů{��.����w�(�0HX��.���hz�ãpX�c̄b3մ�vc��񐣀��s,K��T�'�#�j�2]�}��M	�}
�I���d�"eY��X5����SKV%�Kۋ�p��O�F�aUR�(��r�i���E����ۋ�#8jUS]*5,�H��z=� \�`�n5kl�-qL]��ܲ�2a]�l������M	�0��)���������&��D��{~����VjF���5oAg���f������#D*����.W��� U�z���My^�um�i�0I~kL�7l����JЖ�i��w�hT5 K^���f&�Ԓ�^�v�M�x�~^�%�H3��뗃�#����#sw����2�
�ICX�a�N5��QH���]�a�7��Q��M���5�E%Y(=i�o�Sf��XϐÞ�*^EN���v�%ϡ�,B�,f�K$b�Ї���wCP�ؚ�ND�,��$�5��:�ݱ�-���+�n�EȔ��*�������6;
����)Н���� �q>`k��y,����^���᭕1��KE�.��W�+�m�s�p�.GV"`���%d}!��"�y��d!#F�]'�fR�r�T#\���C<A��/XeC1*�6^��r���[`4
�c�*p���rLX"�����K@M�v5�pV1�h�m*��)a�hާ0��/#�b�gor��r�G�^��q�P�RE���O�e����槲 »��=^�������P9\��G_K�,�r�'=la��N����kK2���x^#�?t�HJ\�/�^#5˥��K�:�͢]��,���9��\z�����6[��vRrs٦�U��e�6�ߩ{����g ����Z���o���0��qi-_0X!=6��_g� �����Z8����R�j_z1/rȜ��'3[Bћ)�tB�� ��Ǚ+Jt��&7��i��?�9jt�d��nN���+=�2�+�׼S&�\��J�Z��W:X}��T";Db�.k�-�j`Y�Adߪ�,�5�`����̨K��U�gOS���~ʒz(�b ;�]c�Oy�eZ2� ��̺lA�]ܣ'���o�75���VPkE�2H3�f(�K�:Fe�*A���k�o|�Up�p��0LrF��j���)/c��攨 [x�`�T�V�#���b���w�fE�9������܆��,�5��-9S�"iŗ~�t@3�g�Yy��$L��du]a|`�-�'�4�Xj���� ]�B��#}R.~�&t#�@o`��M�l�?�A
f[K#����4٥�����T�d��Vq,5M�5
��v�/�.��Bn'o��;ӗ�/Ӣ���gi�x���_X�k5��{s��:�tU	n}sC�bR�8��Wj���Z݉q ��\m�m�LǼ���I8[~;)EQW=�Sz���)��k����D>k��zuto{_u�#�ò�����
���8�C1����c��������f��I����X��dB�gEX�,��I ���IC�@
޼17j�o��?��j٬y���?�EUNɪ+vP��k5�QS���>~�:6�X��ݱ 8��$�cC��d^���mw�2���M��1l�_�����Xf�����������u�s�@v�S'��3�E@O�EG<.���=V~�m�\`ZӅ�Ŵ���0��=w�y�' N�jj�w�xHJfYw!���8�O�d�(�j#<L���2t���:�YS~&�n�	�(�;.�վG4�L��j}�7=ĵ-�	U�����Ò�M��
�RR��6ԴM��\�"��!����t�� �
1_b�؏�>�μ��p�`D�j��q����ۮ�l��q��R��3���[���}����n��L�E���L.������?Q�&$���B����d`DN���[�yhe�
M��E���#�����p|��"b���V	��?���-n��Fm0.8�S?�Ǔ5#~�
	jZͯ����L %�SSj1]�֞�#�%NL�0��$VD]��a�ۨ��6�a��.i2�,��Zh��C���Vjw�M�g
W�Vbb�xq{�|!��%�TA��ۂ�{��B*� �El�hdZE:�ܵ�df>�����dF4�
����!V(�E��(���|�]�/t]TO��Z���Y:�m�TI�2�9`�Xiؓt�j�6��h`�x�E�+K��V�L�mq^ ���:�6R�-ꉣ!�a�Sr'�ą�fX�3c<p�MJ�eM���W��Ƹ�:�%���u����=ҟ%_�K�a������sq~�� d�{F��"O58yke֪���QG_\Ĳ�o�?]%��9��TW=щ3
{�Ҷ�B�xe�'�%��;t��B5$+�uL�y�>�GXD�|kW�N�����\��t5�*�~x,WR�[��ǂ�|�t�s��U��*��ky�v�����DW=kUr���PZy�=D�˝��E�(�g�<O'�.i<ن2���vġ�����ƀِ�U���o�?�Qt� >bK�'g��VQK��?�N��e� c%�A�MP*�SpN.���:O׶�}߮�_n�C�B�wg�"ə/��`�W]�h?E4!�Kn��6�.1L���؅�N��A	z��wQ� P���hC^��@E�P&����P� �'U��'s���@��$�0h�N�w�n$��m{���A?�i����͆^0<�OG�}t�I�Y���r�al<.�Q��A�o���	}����_��l橿���^�K�3N��>`�ۑ�q�0q�,�|����~D��Py�|��zK���5�
�0�Ii���RU��NS?��n�n�M�R�u�xEm�i�J��w�)N�7�.�