XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����D��`]��S�P�"�EN�Oa��u�8z�(/��
��A\dhL�m
$G�sh�yd<fD�G���aɖ$M9\U^쬿$��·ߞ��\w0@��<RL�@~F��(14Wx��b7we��w�1k���ng�u�u���p��Ê<�,�~!#I`d��p�w�k�c���=-|ȐC�wo��,$���
���i�j����P4u��R�ؘk�ȹ�n��-�	E�:� ܢ�焵�̠���-��b�.�Q��1�b����4 hB�F���l�p��Qb�����d������t0)y��l[�kt<y�
@>���S�!���v{�:th
���;����mϪ�>�R�55tm�8�3%Y�:��F�v�'�c�;�/�h,+���h�f\Tf�`H�E��{���|�����tV� i���Q�䬯��I䇓[!i��.5QM���#�'J,<�D����3v�sB�F�9r��"����%H����p1*����P&b�Bg]�D����ϧ�Go9uޅ�O#َ��$�f\��7�}��b`!q0�Z�꼩�݂߫q�������T�};�:_3�������<�����k�Z�R{�9���Q��&-�d\�i0���'�|\��脹>��T���O�0����[�.}����l��F�_ ��!V��P�z�5|��ه~�1�����w��C����!"}��e�ʵ�������������	��J^"�	i��R�R��A5XlxVHYEB    fa00    2480��(mRolE]Ȧ*It����ʸ߬\�e���栯SȀ8�2�]�;��?����A�,;���:��w�4�[�`��ʽ��/�xS;٣�A�.W��QV�2�������R9��y���e����؄����3���d\����L�;���
xQ���2 ���=Q�>ji�%��r�1��o��Ζ�4��,�jG}��b�M!��g�����l�O�@"T�o˷�>���=�D��k}y�G���e����ͮ�#��҇GJ��]&�Uo�@F׺}E�Rzh#�ٰe�_6���t���1�Ȋ����
�}TƑ=v٬���H�7;���*��K@7��C�l����ݝ]�&w{�`�}��7�fQj�v�8&\<�Y�R6f�ɓ߉��ԯ�y�P�6������W%�II�X��3;�;� �)��b�B�II7�2x�eհ����Dl#U(�����+N�'��i���A��׳s6������4T[Xσ"ԟ�����c��q��':�:��������M�^M �8���c��{��FU�� �=��Ȓd�%�f � &��Հy'&�t j���f�&���܌{~��o�b�F���^��C�TP���\(�Ɨ����|`� 1��V�C��7������ �դ�%��KE�?��:�nU6 �Q��ǂ�v���,�:�]3�(`���5h���w���fO��dO����M��G���֒Eᕴ/�Dc1>\!�$���L�y��7��q%>���Q|��7��=�G8[t���o�s�ťN�g�wHR:���H�N?i!��q���T��%� �(U�9ß��s�	5�Y�ڍ��,d�\d���
d���=v�"�rP^:	u����H�u4�Z`_H������
�� ɔ�T�4�.q���������`��Ni.�l�O}h%2�=Q��ʦ��������ݾ��z��.��]L�i|��g�W;�bQq��oP׊�0�oJ�<�KΓ�>y��1��'��?
�.���6�P���Y�RXV�U}����>k���A�i^�1�d�a���n����R������l^Cl�������UR<��9�NP�V�5<kb����L^3��4�G��P�����v{�#������x��:s�s�sJ��8�[C�z�[?�������.t$���7��oM��2��Z�I��Ӧ�x��7�
N�K�q�Xo_www�pm��u���fU;�#�A��:4sa,_�����QRþ��PmE���Iɉ;&8��A��9f���^�ө�2��P�<�)v"VH0�Bv8��2t]A�{\]��F00:�q*@CYP�XbCT����ڡB �%�ƺ�r� aqQ(O�MU�~�g���!�\w�F+�|�i��������y�R�`��Е������#��Ղ���@#d�yK�z	gv р�e]��9G��3�p�}Nl�hO�>�aF'��r��Y;o�I�.�����g��Ú�����{��X덇�絬�6�x�,@Y�N^0��bm�(��T8E��t�b�7�v��m?�U5�x��\���`K�uD<�Ҿ֨Ԛ蠢�D�s�+�$���f��H���My�i8���O��'=�n���ET���}��Ve�=��?p������1������?�@ .>�tW�D�Ww\S�4x���0}R����4z�#_��Dj�+1��>��)��c�~��|Pi�ܕ��.1�ֳ�������e��U�1�����׶ʳR)��<���P�Q �9�lRY����>�vI�sԑM�u;�k��-�i��13 Zn���<_P;�s��x`��W𩦛���^��+��q��6�K�=�2Q�Ň�ͱ��"�Q-�:C�0�l4���X�=W��DY�����6��;w�xxe��D�*������e�~�$T� ����ܔk۽~8��F��z ��X�{0���xiο��/#3��5�E�Rѧ2��{�S�6����������93�����Z��`��|�1��Q��>p�#S!j��绍�_�\�i�.��zG#�a�`ã{ɸ�SY��X����!j��i<�� 6���d>Q�&����8�Hȃ�$1�֯n�wL�*G��9&vW��nJ��K����uG@��<�����ћ5b�{�]3��u���1�Sr�c��`c�8�{�������
������bM}D	j�D�D��Z��!�<a���\x���P,�6�v�+���.�Ԩ�3�q��j֖�3&-vl>�g_�^RF6Q���o�� +���o^��}��g+�O���Ϝ���F�y=��s�z"����ߗW�M�#Gn�	e�C����wz�ʵ����J�D��a�0��붤�πmؽ�S��}͑�6P �1�*h�Yރ�J����'��ōrġvp/�=�8�^�e(��rN��	r���t��
ʈ�\5"��?�o��p�6�FH���v��ǜ���������ſʨ���A=��;�i(�!Y��i/�{<���%`�/�`ʸ��pԌP���?���	��D���\�u��nc��Qv�����a;���~��@���JD`�D��/oS%S��O��љFG��IAc��P����5��nsg6@l�����K��'�jK���q���6���T��E�E�s���A|/2����ۍg�F�X\Pӯ�q�:�.Ƴ�|�ʏ:4OIiޣ����ֻ�D<L���0Ul�b�S�ѵ�2#����ڋu���i�y��Y$D�L�{"<	�Y�H�������4	Z������[!K�-��a�PNo|8�1@"#��~�M�3�������To�t��LQ3�@�l�S+xU6yY�e;4@u�^Mf[��͚�cN|KRO\E+_����gZPJ����2�(\�������'`'Z�?���dk*p&����7#�%��骐�΍�֩_�KG������P���F�8?��c�H|>EXL���!,5f� RIIr6L����3�
�ֆW��ɱ�ϛ���Sl*����7թ/�xL�����$@��p��i�wd��!�;����Ae6�)Ȁm�?��]G�#�'�ʖ�	n��b�bf�����8)�Ą�"�b�8>��H�#�d��b�� ��.��b�Ɗ�+�ÿ�+{��"����ۢ���}J��/��-�灷j�n'����Z����"��T�!��������0�C�K��0uY��/I��D�B����->%�M������}1}��๩K^�2���_��ꩇ&c{�t��?V�ZS��|?��x6zצ�Ժ��� 4��o;D��٢��/��^
��@����5�����_�?_Ek�
�ܸ����.
�'�1�Z�FWp�3������	��Ӎ[�ʸxV3� I�|�����4j�m�B��w�z`��R������T$������5�
�#���P�b��.��ز��F���`�~�N�����9�ޅ�W��m�,*EÅ��'#b��e��B8���f�}Z�Btj6�2�t��/��T�p�l��G��އ�}J�ڵL�TC�&k�/�v&����a�� �?Y�mW=bQ ���E�S����u�e� �O����V���q���g�·�i�ɱYs���[L0�U�lo�L�h^A��ДŦ�k:�����wg*'H�*�E�a߇D�Iʺ�!QϷ�������_�����@p�d��G�h=:Տ��2`�:�,~ž���Hh�#wI<lK�w�Q���ަ����L�W�Z&OW��Gh������/f4�����y��Z�x��Z ��W�M*[܋)Y�O�3��K$�w�9�Ͻe���No�2���� ZU��K�j.�u@�M�^�����Ã�sն�9������h��&Y�A@�H�i��ߗ���\N�GJW�����b���W���ZĘk08�?7R�����K��O��JЪ}:A��$x��<Oo�=wVAe�Ά-�%\�*�����GY2Š��:�����Q~`�k�0d�Lc��ǀD�RnJ�����.L�8�v����� a�e���q�����-i��!�,R%;Ԅ���Yԯz뻐���7��2�;f nK4��5����d�z���-F������L%�*���R�[J�sr[�y�����5��N/�ܧ �Rp�B�����A�+�EU�'�
��v�?����N[e�Nj�u1��S�Ф2��ҧ6b�Hy����X2J4��Ajz ��3�Gӊ܃�璽Pg/���u��iP+��<OU�j�e�_]�*͕ң����vt�%��V���\����B����g�XFj��ο�h
<T�4����PoOS����ſ����A�,�2�|��5��8�X$/A�$�1�f������kϕ�S/mս�����v�>�.�Q�m>��b��ٶap5�����Y~��l�K�p&撪�EFSDv�K��u�)�:��-W��v�_�ϔ"�����E��ވИ�&�j�P�������~ ��0�0�c�Bdw�#�pbII���N��,��2	#ݭ�f:{�"v4���5MKf��nP���Țͼ|��!��猘h�=��@�@��6����V��/���1�<��@�ue���t��~���ꔰ��qo�G�ԣ���rrO�2U����da�ܻb�엍�Љ�LI/���c�<��^�U��л�vx\�pJ48�.�t���P�]��T�Pm6�� h(`�V	mQ^@^Ր�TU;�r�:Q�AI�ϯ�f���J-F�h��S�|�{SOvyȿxP,�B�X���N]K@��k��r��0�ָ�ѕ�6㶺`�m�N8;�y9��N���$Qe��j�9�2��#�0�Sy�f@���G��+���-YTxٕ�l�Γ-������gK�MW��0c�D�MоWK��1�u{��~%wK�IT�qY}���=sU)��Ԫ��F�)�D�`����N��T��POt�^0�o�#�xL��|q��W0>D��f8�J�y>�]^cÔ�P��A�ϴ�/�V����7��9ϴ���+�P2��o�!�����vMvl�x�i�:�%V�೺zkCLfO��3�2:v��L�-��~�#� �U����Pi��l��]?��^Ҟ��?�[#8�%� �Dts����U]gi�/�+��]����#B���p�^�����+��]�H5��ޒ���lO/�6���#B�z�'�b�
<���ă�v�V ػ�����o��Z��w��π��gps`��(0,��a%�抮&�(���
 ��OԀ%<c��N m��?�&zh�v8bPKb��N�>��NbJ�ܼS�R�������9�0Y�.��\��}�|^r��S'?Q����a��vXS
7|��q��X��&�!�i\�c�
S�����}#�Ѷql�9K5�@ȴ����ȓU1����uXX�g#������7T~�i]�
(�PO��<BP�P*�Z?go��¡Di��	9`�ad_�2�˳ �E06۷�ub2jtI.j�D�OR���f .{I��ʊ�M�T��߆�J`����ѝ�b�'OM���}-�bŚJ����'��U��y�@Α��Iu<#-��8!0Jc��*=ԅP �U��l�)��g|d^�L�T�f9�:�O��ab��l��,�%s.��i����^�o"b/I�IH2���]���r���;̂����b�b���$����6f��#"8��*�`=�d��yP�m�8X���ⷠ�9H�ض�^�K쭻.g��O��*��9�޿,�
K��6����|"��)�!�Y��?�t��|ׂd� ��*Ԇ�Y.�S#/��AԱpmX>GD�5�-�yތ���rn�k�3/���LCo�p��j���������[�:���2Uh�@��{�*��,�Y�Q��Ca�
�c?-�y69C��F�"�����9�P_{2p��^�J�g�w8�u�����۴�"� ��W�:H��`�
��K��ɨ"�L�T�ܘً��7�F�;�r�Iׁ�~��~yR4�o��(B����4j����Ԛz1��IB����X?6�'�cf{� (�vg�l�����{c`\�O)3�ˑ��+A4V�aZ2���V%��U��D��C�ر<��`� �H�f\�r*���a�KebP�Υ�<����$rg��!��(W�y�������Tq{�塞��>t`ѻ�3�|.�QK�1�%O���VE��p�N;�����l�^?
�6C�W�)%��CJ9e��j%qҼ�e+��-�R�.�lB�r0�g�z2��.y#������'�E�5?E����������L��2؎w��ϭndR����\�x�2e�;C�!����;��T�"��K�T&��$4#��c���t2���M�|Mf�Ͻ��̰��Lq��Y��D����O�.�B��+��#�a�Y�U+��č��n�}��=��H�!��/���S��p�{�JKt��U�
��N��H����]E����\ڹ.��چ�F��L�6w�n�UK5��&��=�"��D�þ ̒(#��BP����v}LQHh�4���ծ�]�P2�i 5w�ɑ,,܋�a�#��;�S^PR�Oׄ�M8�%�)@�.�4�7��}�[�W���*y9�(,���*�[�
]-��*��a14X����_G2�w������������!I�=�?+��'�[�d.0�e��F�/�"����gW�Ѱ���!4;�ːߴ�{�$��9\'*c��1Ih19�s��KdX'�k�ô/G�2e%�ՙ��b/���2I'nl�7T����,1�.ʷ�R�V��T^p>��Kl2�]7�e��a)�zx�-{C���>,= ���}��ؽ�j�H�box1�5��b�Xl�:խ�{�c.�Լ�q�B����6��O�X�\��!V�\�o�;ӥ�s aT��@��~@-
�O�)���5�^�dc.-���>Q�#�����go^�(���ɐݾ�%Æ�o�c	����a4��W� ��� y���K�X �Z�,-�\wFj0?�F>�l��#�F��/]�����Cu���Ӽ�oΩ�&���ޞ5dw ���o�z��'�q�ц�ѳq�oW�ʋ����{��6�t:��O���G@&��e8c����ވV���m-��ny$ߪ^R&͔�}U�"����;I�`,�Sțܢ��!��|�xR ��8}�Y�t��mLcʭ�B�Y�Έ[���{3�w�f�(bkin�6\d�6�l8o�^��xK�4
�ޕ?���M��t����V:j��κ���X&��\�򷬓;�v��.�:�r�У�g�$JeL��(����TW��AO��jM��y��'�O�4K�o߀��[T9�Ok�ߡ�=b����$��J\�6�#���_��qȂ[l/<�K�6��pc�?�|���қ�],�����#�]����i Q�+)0%�8�ڱ��;I5�`�sF�h�v���8�N�w>6&�&�٭�mt�`����M�����CFeVW�C�6�z��YU���QN�(^���Y��Ԉ������@�x�Ż��[�����ػ<ZF��W����r��TS�}f��^�;�!�{��@dz0.�E7X�j���70o>#�v%�~�CKbM��˾�Y���7l�tfp���[(���'�����}����3g~vK�'�b���K�5�:��P��u�0�#���a�����DG�U6� W�� !�k���S�*��U�e�0���b�}����B��/c׿J5����O���S�I2qތA8L=m�	�UD罷��$��Xߜ�!�I(�8v�r��X4sf��]�~���ëEYQ*�J��w"9H^�u[z��3u�*꼨?�a���F�v���j]y
���z�H�嗖Z͌DO���������[-Xz
��'Dh/����G�=[���E�T�/�X|�o������W���&*:ƶtt@��6���8'&��;tP����`<���&@�t'�+����o���)f��B�;���a�o���<(\�_}����k�J���}���C��u�@�	p�~�@�Q�k��Wn�$G[�8�1���K���Xw2"�Tq��']�R����)1���H�Us��,�@uC�'\W&�+�f4���( \B�h����ȗi�T�G͝V�����خ��R|�ZO�HT��MY|w�T7Ns��ϐ�~�-;u���2�qR+��	h��Ը�4����m����G�ޝ�Uʺ���O���l��5/Prw���[�e���傠K���;�t�씕�!�w�W��>Cp`.y�Hl�
����I�bI��X��4<�cWBgP�7}����?�����(~Қ�3�R���,{zr�Z� �5��=�����8KW�p��8|�F̹'D�M���������ZK�P�NR���eG���3�I�v�AK�I�7�5=�4�^t��Z�lQW��KmW����ˁ�~�$f�i��q��jJUVƤ�y��1 �cԉ�a�5ަ��R�I\S�T��:�:�I�d�1�8=ρ��`$#>������ay
>BW��r����ʢ0��*ӡ�?����+�e�h:�×3Y���n�1S/Jx&y!X���/��,[4���İ8�p�����,e������Y�C4�ϋ��f�5�&ըe��O�UU<T�'Ǳȕ�6��kXN��ܧCx.�`i��v�S�R��O��w퉐��Ɋ�f :�ދ`_]�	��A�<���ʛz��bH�%��N��X�~���*6�e�$�v=T��A�[�����>Ϟ �7��8�Ǎ�ٺiT��F�7��z��k����4�Y`4=��{�� Cl���`�l��c����*�i���veS"�R�q,������+tcRy�}h�_�r�@5� ��Ͷ���iٖp0�l�A�Ka�:���0��Ֆ�7(�
E�v���A��$� 0�F(�?Z�&ƨtX�e���Q�gwC��Ҏf��R��#�&�t�(0��]�iK8��)�G쏬�ٷ�ru�^GI����
o$?�%H�T��N7��oTPl�I垯�LT�.�AK<s�P�d0�L��ˀ���N�`t�4;�{l5ͯ'��7�?e��W3 kn��]9���d��?4i�XlxVHYEB    964e    1150���+v$KVx�x�wҟ�j�Ք���E�t�g���F����2��#�m�1��i�w$5�H�Qѣ����K�z�+�L�|,�Y��Cz�Ǐ;?��������XͣG��ۖ+q�/� Ѫ�Zx�M��&r���v֩�*�VF��cl$Ֆ;tfй��~6�Ȉ[o�tb%��[���e�)��\��`b��M
��Խ~��$�w��dE�:f2@�FL���]��V�v���[�	D��'�}��>}Q����!�rV��"�4��	=��T#�W���X0�ʧ��*���ׯQ�_e�aV.�\��&��^@S���)U�U�� �͒<=��Oa-����Xj��R��c��B��E�#3��Zf�IBuؗi[����r��@%��x(qx��%M�<"'Jf�6��� /6�}q^�j����d��s��W	gezU_��Խ�k.Y����� 	0�	*�J�"%L��DyW�)��t��1�B�\8hҚ�z�c��������A#�Q��;������� ��҆��m?��ϔ&����ez���3>����ZrG~`?��:=l}?�K���N����vvI���%�H�Q�=��)��5�sy���^����Ydl��_����w��z���(�S���7�ȦT���V�?%�[p�h��4.�FB��E\ �ڇ"4LN�)����a23���T�k�y������c4
�P\-�+*�HءZ6Ij���W\����0''�I�˽��(-�ER�|	yG���.X:H2)�k{��!Ad�dB�u�B=�Q�2�=7�;f0��-~$W�w��w����-Ye�T�l?r"r��&|5�w���׊�5Rv��0a���
N�B6�;��+S�T�����M��A�`|��c��t{⼓�}G��9�A�[p�P��w�=��`�o��/��$�c�u	!PuL�5��(�*%T�̻Қ��#h��%]�` ��kr�9��qt���d��)w%0Ī�rỴ��L���5�▀L�bM6)��P�m�ېӆ3����<��у�>��x�E��>÷�byo�l��`8֡�o�g����%E'T��|�v�J���.R6�t��� �rJҗ=�Y��H/�X`�6�}n�r-3Mp����c$����ɥA �,��,̐�i��}�ĩ��BD$�+q,;����gʐ��N�>�G�E�mم>sn�ԗI�T$~��d�'�5j�J��l��ՆW�0�a�� %|ټEM]St���-}�Ru1�Rr�W>7�Uʵ	n�i�^���Q�μ��g��q�������V�F�V�zv��#e��E����]�R�P���{W�j��[_��#������\"x�7N.+Qdƿ�(9���8�^B�7bc*�`[Xu��_����w�V2c�J����	�h]�ح*w�D/�$!�����)��#�ɛ�5�vѓ�{ MP��­�� �y�<��G��YG	Ih�l���o�s�՛�d��G���>З��1�sm;]�M+���Ž�ң_yB���� ���m��<���!+�u[�%/ ��9m��eq,kD6�sX�O�KSf"��:͓�A#�� �]������,W�%��L���E�[�p��3��#Hs�no�W�mB�i.�ŶԽ�;���;B�|���.h0�nN�O[�Ҧ���,��7,��@ѕ���\;b�3N��l��1�z���(����-����8!(�e�ա�g��Y��e���M#�+�W!�,�@���Ó���C�����@�kQ%�;ޞ���u�6��>X��W����Z0�m'sq����4�>��R��;2β��d�Ng��-:l;?����|���Hԑ	�<���Js	���9����3%S�?�$1�J�*9.���?�b>Q�ɂ㳖+�w�H�cyq�O�Hn+��R����V8�b���M��T�<�F�ʍ^�$Qk�
1QN�9W��/��7�RZ�����b�M�/΄�$��I��W���sƃi(��\�3&��)P^0��pʦ�[��1�U�H��#ꄭ�@َd�&��;���\��c���$釱p����2�D��oh�U���H&���~Ԏ�ᡫW��{� �Pِ$qǬO3f����lۈ?��i9���Vj�\��P `��'Gi�7�����e��ùޤ�:dt�����N�Wy� ����m��=k�\�S�P2	$�S��P�XC�C�����K�ʛ��j�G�<���/6P�d"A�5ֱ�Ȇ��f�C>#�ǈse8bҫ�70쩳�����u�<+EyV}�RQ�X26��q;Em(��<!;]����$�'�r2h�����7��^-�c�uL�X�:��}ńɾ�5�x)���i�!|�b?�	��]pw�y�0�F���'�P;��۟��x����+_r,�z�/˕�1+-�Ϥ�c����bK&�`���9q h��^��!*�`��n	:�w�}�� ��	�����|\r�F�=����#����E�@Uj%�J�z�p~��54~-!�^�T�T�G���g�к���@J�n*��R��\;� �c�̹�,�8dwF[k0m�AC�4۰�B�xO�=��&"��S�\s��E9���.4PH��zY�8T�@� UJ|�}�eX�c4�1n������ݪ�q�ǖ%tȩ}�Ѧ���z��bv[����.mf1�s^��Ԕ�v]��Ŋ1�F�~S��·x�rQ׉���|7M�.k�~�v�����j7OS�$��`S�U�c�ew�NS�l+����Ⱦ:��`��>X)�8XCV��%Y	+�Լu��~�����$h�1�T)�q��YX�m�̪$��>����T_Z��q5����m��vd
�=3p�Q��A)\�D�V��Qqa�VTuIIOe�i8v�!9Wś��ܶ�-��H1ں3twO)z�	���]�~Ѳy	3�?���	E �;p(��}���j�'>{�(j��G�ʧv�oȞǹ��h�Y�C�"N���NS�ñA���:���U��Y��0����$w�������o�q˱ޙ�����.!���EIM1��=rUF�����b/��ݤ��h�Ǉ-����[	�D��C҈/�;���k��A�����R���)<�0F��d$�����E��f�9�_���uD
@��Qx�D ���Ø�{����2Ґ�:`VEFcE���vi`�0�`�M����,ѡWq�j��/n��?%���U$
�����u���@`��`��i�0v4��4f�}�,tә��p�GD2ʷ����lY,����;�g�f��k	y��������v�\��[�ŻZ��Dܝ�-+���q�lsO!��u/�����ö��[)���|܃��,U-0?H�qD������R ����� X @B�� ���xv�OM��KN(,gF����Y+6=<A�P_�(>a7H[׷��h���V�w�1^@,��ޅ���YC4��C�n�;�lFy����8��o�C�����I�T�1�46�rY��/�Z	��B)Fr��X�r>��œp�g�^'���f��<y�ed��!�;��~�P�D���
�?D9�I��ʡ��C��)6�9�}n�82�W�i���l��&W�t�R�f&J���B��7� )�vWV�6�J܈��[0 jC[�n����R�8G��SE[;�7b-x�ﰩO)�rvNjfJѻm���F�����]��9=95�OS�&�!ִ�k2�Z�3�6c*;��W+|��e��沼y��D�6��Y���g-]4<�LU�j%�3�6B��#�X�P{�W�Q�c�~`��i��'��]��ᇟރ�e�z��tX]���^5.��'�bd�Ɨ�ĝq��_�}�t�4�QG�!w�k���.�j�M����V@��h�S��h@�h`$��1����nuqt��m�L�v>GSҫ]i0���q��!%��Ty�K��ω�bbg|��0v
�p�'�ࣞ�!�=��a�s��oK�/:���t�Zy�>h� z�����@Y�Q�0���H���Q,�k�Պg�Tt�z�z���|��o��d`�b�q��)Z)�Ȯ��h�y�c2 �Ň�3Tc�Z��*����͘�"#�
�.7���N���z�hX�6_��
8QvB�ۨ�{�`(U�>V�b�J���0�n�E������C��k'F:��y4�7Y����݁��%�܇�&>�0ɸq/����.���y�yeq�U0�YS��)
�w���up��=���x�H���F���{dl~�W�L<un����6ZQ���n�yڦ���p��[�ʟ�@eXïulm�����>P���-Y�wY�a