XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��İ*߳ZJ�I�{���l��g�ǅ��]�~���P��f0/}?t�=l���l����gJ{�^@o룳�w�b��9���;��478�	cPP����&Rΰ�A�a�o��{� �G�j��sO*/m��atQ-hlߺ�rw	�3$���9�����р=-�_wV2��#��1�� <�z7�`�0���g�R��6�V uˡ9�v�X�NA	*X��'�>;n쌇D�����{��Ͼ�lu�L�C���W`�Kz��6[C����>��P�
E�Fz�!�>HW�������S�$���fI��0�v(�mz�?%
��
e�fGZG����;��u�+Љ����$r�{���` �.Q �<Q��:��r��������#��@U�&Ӗ˯~c&���8��J�/K2%���7�H�)����S�ީ%�_q�N�~�����/n�?����������/ϱ���U&��ꊖ\m���-&1
��)��G�&��W���0$�K����XJ�v����Q9��Q{(�e%��;�E�腟�;)E�V�MԺ�5��X!G�w�$��;Wihת��пk.]M��z�-�@�z�r���␶���t��vP�-�o��+%�5%�b�`gN�����h{_��gV)�;X�,��&����íw��U6v%������W�j=6�w1}ż���p�k`�8.af�3s'LjI߆=~n�ĕ,�-��V/^a����+��d�nS�dj/IXlxVHYEB    7ebd    13704�(�ଉpwh����:��Lz�!��/��+9 "I�X���b�`�~N����jC�)%'�y8�r����#��2(�j�4�����>\J�?A`��>����UH?�>%��))ak�����!l�Y��G!�|σ��e[˗aw���$aH(NQ��DA|n��2�����2�'��t��_)C��HhS����eTI��̬S�OP�i�8�9�W���qO]JlvB)���ĸ�F�D^қ�U�%�g��!t�d��s�I��{�����pى�z�Z7i�.�b�@���O�"g͖�7,�~�A�l�\�ґsV;�������0u���*3q�M���Π�<U��87�(a�ʻMmx�;{q�F�,��	�DI5M�ҙ���
ddF��7�NtˑP��[x޺=�1�H�x��>�rb&�-5xX%��?)�h��nb�F�c���ʂ=�s�)�]��zR������z?U��%^Ȩ�U�Ҝ����Ν\8��V{"�[j%EZ����h��&����������F��.t[�ݼ����mA�|��br�����U+�T�]�&�����;M#� Q�A����˽�VYt�J��O1r�xۏr������x��`����:�63��VJ�0~��0Ք�vط�;�	��k0�*���Ӟ��(���o+��s`[���&�X
i�y�9(��w�	����fy�H���[� �w�ܪ�˄��\�*Aq��AUn*.˧�1���@D�+Vh�ו�U�s��W�eU�&G�+����2E�uc���Q��eϱ�ې42��k�4��ߥ�� ������?�<(�҃GO�H�A#f���I�埂ʨ���d��vA�	$Ǯ����]�QC��M��k��"����GO9��=�|��{YX˥E�e0�RsLW�Ț�.2�_�K#E0E'��_�u׎�e�i�E5�d�XO�gTz�BB3�VoY��T) ��W��c�^��r���3�
��CB* tc��U,�-�N�2֥a�V��������5��2k���7ˈ7n��3Ynn�,���]��3��^CYΦ!Q
�]�:=Ƹ{��˦B�;.b('�A���s���|��#��r&}��U��oN��3�)d�R�� j���A$��s8I<�u���<�C/�u5��<�n�&�����R|R�ٔ�AqT����ˉ�����u�4=
S��)�P�d�<��'%7K��o�F�Y���B���Ϥq4jj��@K^%"�޻��HȤV�2^y�q=*h� {'�k>*a&p��N�W���d�)��M����\${j���֬e�n��z9[���P������8P����j3���`��)�O����IjR3���co�/VT3�/�A�����OS܎t������1��	�(�R����&75S%dH�#�ɛ�ͽ[I�3T����H(�
ѡH�ʩ�to������׎;�l��3T�S6��0��^�E�\���?]�bx�Tx@~����u�Z�أ�!4B'[l�]7×»S�;*ׅŰ���8�����B�r�<����HH���n��NKϬ���S0%P(�W�FxP��r��?�<\0���ܐ���K����눴ō�Zx���@BE�9jn"yj�?g`С�~���G�;�	�N<3|xK$j�+9�7���'y�P�	�k(��@�%N��ؤޫ#��^��[x��UⓈ�uX�y���R�����~Y�f˃M�K��R<�D\�I�φ�2��>�KXʃt����Is<���8
�V��!3Je��j�)�XWG�J��~�G��+� H�&(�ݚlRk�\�.�H��'�Nax���-(hd��[2��M��C�}�|��TVŃ	�wP�&8�?憩�����$�"Gl�'t�t���Z�P2���1��|��F[,
"�m��F�}�*z�	�_��Ȑ_��wC��P�H��iD���h�s�Hz��El��59�먑�H%!�rG��UNq9�́k��,��{��|���d�����uś�Q�EQ"��hEK�R-�U�H�w��5%��U����w ��r��h�%���C>��'Yul6,p�֭�x���w�.�1E�Ճ Yt2D�~�>'�ۊ��7T�6�d�L-��iΗDh.�Dh��qU�-�^���_�sP%N�۝u{���,���@C�r+ք��������j��5�a��r���GH��N�P��� $o/d�c��2,l��!�ӑ{l����,��}�݁�M��
��@��� �%Q��Mu�L��X,k��5����R�(� �kr�A�]U����>s�H\@Ӵ~&f
�V(6����	۶��F�q��k��Do~zm����-���$f$�)�9!��E?m]�ǰc3�H ��o��N���C�a�l7�#�2>(��(�t�����UM2���9-�[�^u�f�w�^V��o[�}�{��1����D^y�% ��z�ű��D�ds��f֠�R<0�>J�1�O�8�.�-'��.���	�l�&�`�]8���-85#?/2�2���ma��x J�{T��nካ�N.����*���Kv~��Dh<"۩ґШlg]d+�عvI����v��u�L�Ie�5!�mr�,�ҩS�J��4y��\�R�{��h1fܵ([Q�
�J�?:�6q0��,N�W�Z��U�I�PK[BY��쁠MÌg�'�tPL^��$���c4�R�z��X팕�K���]׻��V��o�(��J�9�u���Ɋ�́f�Q���\��ܖؙ�EБ7���KX�o�P���v���;t"��U`̬���^1 �D��6��3ښT�
ɐ�_����^�(��Ɔ�A�{JX
D�csX,p�ZW�SA��w���$���^�8
B	��6L�]�.��E��#�?&��Qʱ�sm�U��;�2M��͛��O�?���b�cM�g���q�@�t���&wi!n�����?!a�,��z�4Ѧ�K�n�oV�Te�91������[5Ɋ�|�ܧD-nn42i��'#��� /�����ؓ�v/>玛^�IE�ֈw��EJnVZ�0�꿧`�2������NVx�6���~�H|
��f;�f4��À��Op&�s�%�~ʣ�B]EQ�i����� F^vf�?��w��_ZZ�]�hWIV)�����a)rsn_��N��[U"&��b��� [uZ(S+=�ɸ|J��Ƿ.����m�)S;�FD	av�%�X9�a�y)3v�_I��N���L\Q�L')HQű�v�������%�S�v�����(�v,�@V�RXm��a�s��q�f��(�*���1�� �! ���/���#�/�"<r�y"&��8��R�G���9arm,�.?2��@fk@r	�_��>�H�0=����Ĳ���$��881��|�:V� �7�6=}RXah�BU|#�_r�i|M�z���  ��2V�A{�?��v{�]|O�o��3��֗B&�Z�ڡ���<�J9�q`��Ǽc_��/�	�@N?�����O����S��[S��M@�n��D?���Ta��W�P�$���+mϢ��fsr(���h8�PB��=C���fH�už/q��QjJ��r�cBr@��UD�_,�|e����8��\��'�ܙ�8\F���%(�n��I�r濾K��qC������M������M	�wVz��*A�0DC#���;��H#SdԀ��b}ڛ������z�������ȷ��b!��h��D?��A��VӼ7���^��|u�F��#��J��%@��P�}%��$��q��5���m�����ц�yKT�<��Wlx,
�8��.8(�m4O�a�4���`6�;���'���:�]z�x/�֢�����I���h���5��^��+�In�؄U�_L2�5_�B¤c\��<����9*N�q#�D�f<�y^ۄ��^=ě���@��Cވl��>!���ϴ�O��B�0 'V�w����yU�SQr�uv��I��ְ��Ӓ�"�\�n8:%{Exj�6��lC)]JJ��D�+��3�����PE�-&�!b�æ
�7�����K�a��/�t��C�I�^�0I̢<�o�t$�R� �Sl��U_VM�S ��4]>,��)Хy�~}����x��V.�+���:����65-6���
|嶝�y*�M���=3�O/D��M��C�,þ�'웫g��]߿[�xU�%`�*ѷ%o�|����Ġ?!�#X ��A�~�+�V��`$4M'��4ԩS&��S ����y�\@��7"k�%.F�r��ƶ�;��d�*M@�<��x֪%d�b�a�)}!/�0��� �\����>󾎥��!cq?�(�D�Dl�^���+q�@�q������8��M��� ��V�5а-�͒�)��v�i����]t.)%H�r,�>����W���.�Q�����߬��U����u�I�Y���z�V�����ƈ�0�3��yq&�n�w�J���O)�C�{Km�Yŏ�U|Љ	K����s%J��
# �;H��Z���7��/���w���BKVch)-�M�f]$�f��I��e�ՠֻ���w�+!`'�H�TVk�3���v��'�}��.�A$��Dv��X���Q~(s�qH�_���L�Hy悴ZY��<]�=ۺ��S<�;SJ)�u���˫P���9�7-ErW���I��Ȫ�����LT
��:����K^o�����{n�����7�~x�Đ$?5�d�����p�7I_j´���HϽ���4y�?��I7�MO�ɔ/�xp @ǖ�6K߭^hky��s����ax$�����l[�u1����8����2�je/�Q�x���=�.g�ӕ��Jx3��f��^[��