XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���V�}
�%�EFYt ��h~e��6����\���V]���u�һD7}������?}�.�]��#�T �o螣n��N�Јx���Fܥh�6I;�i�n�P��"7�|����ZU��w�خ���	��ɦLο��Y��:td���	����%��qU�$�P����d��u�Xg���?����CL�a�?�/�b6urX���Z-(�4ٌzY����0�Sm�Al%�i�~g����&��豑�E٤��h��+���%��)O6�*ϡ�_��Da����pNy��٨�� �Ǚ�[X�=)+�ڔ1���j�/��y���{y)R��R"&o*Z��4�$}! [�����3��M�-p��(i/�]t�T�>ŦǾ �#N��m@��TC�8�T���e�Z�#��!�Zќ��}�F��N�VY��ek����R�x3^�SqL6Ŧ`����� �b'�ax
�������Z�.���	Z�d!l^1��?�I���T|`�f)�@�?�0�Yy�����X��`�&t_��uzG/3	6�i���MX��ŢS��gm@��넾���0�Yf��)z#�4�J�(P!y��F��.|��ЙQ��_�{C��c|b.0Jaп��@�e��Ac��Ԋ&��^�w/��U
ڻ��X�HME����+���,�ׇY�te��c�F;PA�u��R�Ԣ���s*�M�nC�7�m1ͻ�T����j�{[���;n9�9Y8���'	�����D��G�}r�\2�1����h�^��U%����XlxVHYEB    fa00    1f80�"k�^-pk�ߎ���!qo�M��#ӊ�'ԋ�iN1I�G��\[s���Uͼ
��.��u��<	����<�hڝ�O�~�\6��^��u<7��eTv~BI&��cz����(I��ۋ2"�ǻ\f#������q�G'�*�1v�e���[ ,-d��6u�!�>x�L�@i�.0җ��!X�F�t�����*L�c�KQ�&�,�a���x9gz��cNhO�"�/���\nZ���"�$�v�����Kǉ��f4��s�@e���i�,C�&��	+ц-�%�Sw�B���W���q�a�>�$��-�	�O�A��8�,e�Dm<���v`я��&8�Z����Y+�/�-��?k��K��V^1H�P��U<�28����eO'�,7Қ�7)	��7C���`)+ �;Am�V���Ө*����n�̲��V�]h#�8��E$��gc3���s��3�-#�W�'c {�bú/�T�G>���O+���v��bbٹ�d��#5qз.�y}^V����C�=W���4r�ZP�����x~�m���f�O�P r<�Ԍ�.�!��RAGR�P]� /�b��"1GT��kL�%�c�2����6��UUs:9���O�����.S� p
�E���D㰦R�4��:.�!�
x��џ�-%�[-
��&��7=�,�i�-�w*�[�^]&��,�Pjp�n���S�?�Io�������ʞbC�N�N1T)2��r!E�����ܘ���b)��f��<�f{P/�,d~�O|���M[met<���������A?�2AHQu���oy�?{������?p��g��ٮ��,��3�����g�bٞ.���:@��m�{��/�)!0"8I���z�M�U ���%� Vy�}�`׵�j����� �]k���c��4ȭ�Ն�:@�,��F3�[ޠ��`��t�쯫?�fI
u^t���m���`=�_J�ŗ,$u���x^�!7MRM}�2#�F�M�������e��7�����7IQ�#>o�/���(�s�M�n����$��s��X�3�Y�!���W�k�����H���JFJ��YF8yv��<ۓ[fG�nm��^Մ^���a�"|����f��_X�x�r'|�PX$��"\�3�����D|}�/(sN��CR,�m*l�8� �Ҽ1$4M�+�L���`�*g��q\v�����������$���m�
�w�l=L6��DTcWG��yǶ�ݮ(�K4����F	�Gݪ�������U� c`��#�0:_�Ҕ�m�g��(�	�) �58[�c��L2�Ux�j��糍��u\+婫�Qa7�tҋc������ǰ���#��<�KP08�NPvG$N�׿��&^O��a��e��;���OSmM�����܌�7�R���� (F;[-���k4PnǪ�~��S���汆����[ڕ�s�L�h#�Yu�=`˻�Sӈ:Ӂ�X��&3��h�CX�~��
��%SF�]����ɂ�`��M���"eSV�)�o�p�7U\�	����z��g]t-ڄ���2���ua��ͽNa��}[����Kk87.�A��\��zLrᖌX[$��\~]c�|j��K��#��0g���AǶ�a'gmZ�m/I���̐xy&H���&ѫ�&a�ZY�R�b� Y���~}'�+H;D�p{<$V���.^�=Z�V�C�iz����#1�io�P:Ė�TNt����K��6Njv�ҟ&�W�AX�(p�珤�bp��^��O;4�T'���]�ږ١�y���J.���*5�Y�,��DO�=�=��኷��ir�����Z>�8&Nu���ne�����C%]�p��I��E�/��LE6��O�$���?���|:�*ry����(f~Cb�GcF��(��{���Ѿ۞9B�y�hˑ"�H]�vzu(ʕ@��4.��/b�o�q��tH����̓N\�&�i�=@0��w��,Lw���b���ㄥ�U�!�u��v	ND#h!�p7�9��^�~&��'�b�Q���{�s�&e?U冰�8<��/e��O?Y0wc<��"�5Ôr<����G�-��Vs����:v�����-���FT.���\����(T�����ùX �2q����K���G�x����0���iV��H]Xm?t�,����7�Y�]�1��xf�K� g���5��E���IM�U1�8-���T{���w�r�j����_�w���OºY�\�@N�n�;u������U��0"��3�7�?O8��NT""���$ÚR�6Kܘ�1�M������OG ���"4�Q�O��Gz�K�p�z����-\(0�69�x��_[�Y����H1Q���s��z�#г]�8Y��U�¦ם���VE�ًb)�ߺ��k�����˜N���P/�϶
{�4���l:z��:�������F�<4.�£˳^����_�b�r�%2�w�&�޺2�6#��+m����7��<H(?14�y���9�o����	�Զ�`�l��;	���I��L����;�֙�fL��N���ì�j���	�jY]�-?���W��<��K�#m.���D�"1�&��f溷M"�������1�#f�W��7�?�O���b�qGR�1-�	<�}��-�"��'�э4�R���s��o����f���[a��b�'8�04I��}+�h��Yo�������
ηNĥZztw��o�G�~s�^���A��3����kfx/��q +���d����·uB(A0��)�d�.Γr�l�%�T`�l���9"Td��O+[acfW��ۃ:����V�?����ĪE�ٯ�rF�m%�_˳R#GG�]���Fj)a�h_|��J�c�,�5�<�UCV�`��0+��B2ϥ��|�U6	5S.�� �_s�}�[ǹ�~���\ە�(�L�<�3�=0z�*���#M�iO1�UM�f'�CL=?���#���ܚ
�MҌ�������_C6Ό[m��y�������r���}�v�ᆾ?��~[�fm��qra�s��"�|��Bk��A�P8b�U��������-����u���Az)C�������������˰ e���zuU��4X<WI�Z�F�Yf�艤�>��
@P�$���8!n��͖w0z1�!Q�v���O���B~�&�F������G�p5�'~"�J�Tlz(�����|�8M�4���N��UYc�=3���R���8��ŷ�C�zn� ���{��E��#����.��Ϻ|�m�_����3�f�Ӂ�`�^p���EX��;��@��Q%*����cq&��lk�
���q�w��Ws�A����A�t�>��)L�,()����ʍ%��d==����x6@Epz':����*��� ^�;ܠ5�r|�����z3!u�s���4�2��x�I��|�+���?5�Q��>`�t��[O�]a��!�D��X8�|
�ђó�T.凼tm<Rdc��I��i'ua��t�uT���b."��~\	+� ��~h�p�m&�2�U�O�vq��"�{�g
�������gs�`�/�h��8�G�ZdM���+�<�W�+�m�/KS�X3��)>�7Q��g2�GV�}���(K�*�w�1��%���S������iֲ�,*C5T4�d��1�K0��it�����?��j���1w ���[��c,/{���S3*h?SUNA&��X�+iC"M���"l�˖����=ɮPWTX���e.� "��\�����2_�v��4�d��!R�~���Sut�hv,�Q*��>�����>՚�S-������ �ɞl6����n��H��K��[>���B�[`f�n��YX�p�}�g�����B4����-U�i[��Is�F_�y4�O��C�P���
+~�'ȝOIu�ʊ/,\ݾ0�gaz��SB{>�zf��[n�kVB=0*̛í��6D'[��U�Q �}���*f.S�k�:��Žh�~&l���DiV%2��5�B7�p�<���2�D,��a� u�⚉�D�N�G@,W�T����	�p�ю��5'O�֕��A$��2���^��*�,U������-�Ջ��ac�b���8��/��~�3��4t�?��M\�i7�\p8�G��Hh��4�w��{l�Eހ#�h�'�^��)��o�E@���+h0��}cU����Pt T|��!���N��oTSm ���%}v1�� �Q��&ɪSzhT�*�%���<Fmr��B����E���;�Lt*tc,桙r�3�Ը��:F�W�x��Ռ��9f�ʖ����J�u��>W*�0dNs�-!�kE���ί�����ñ�e�ꎖ*�:7x],厹Y�H�̶�!��RC���%.�{���J*M�k���xR��`�@�]�K��C�,�AO$aY�����S|Y�s�Ɩ����tdf�.r�PŮ��x(i�_�^>�R5�����7K=c��̂�Y֠�K��q�������9�S�	%��g����"��P����o�*A���_JZx���TPVj+����/q?�y����k\vҥ���Sxۣ-����ħ��p{ä��;��j��T{�C�Z�F�?��E�9R}T�4S\��'$U$��F0fg��j0��'���u6���>(�b`m�(��\�,�Xi��y�5�F��'H���m�K��dU��f��cn��d�zx.*��8��A}0�Yʳ�Z�ޭ�:��Z���b�,>�&�0e�x�}�`��mț�\�3�S,����;�#F}[�a *�:N>1N��
����+3��V>�iAꙿ�Fv�	B�C_��H%I�RX���������KF)�xw��b?7b��H�a��}�6O�u~�����×_$��ߦ��+����^��^Ӎw#���W�	�N��s�Syy&��RgE�-�nQ����	i��p��K��>�#Y��(Z'��S塪P�:��:����1ly�y�������8H����;���þo�
�
��_[r}êZI�� &9��3Fy�^-憊��~-z����w���b�l'/��E�w�>��zJ2�=�/Z�X��6Wg+�IS�M z痙m�чs�'�U�i#Ȩ�c�AlIA���)6-w@�L�X�����e|��H���ғ���'�(	�ro��]
 �87J�&�b�iSp�_�&��C�.M�}�ΐZDf1	�|j���� �J�����Wo�âb��"K����	Y�ܭ��0��}���]a���JsԷ��6j*I.�z��[�v��a�������2�N eY7���D�}�!�[5$]�3��V�PYu�5�}�|O��|�B&��ny����+:�ph�	���m���GO�0��i\g�ߙ>O^펫8�Z�?�%��^{5�&�p�r��r�yd�w��py#����_���;Oo��ʳE��ބW��/W	*���ruWC!:�	����������w1m�~���_�6��u�9����vx�n pm�fY����w���Z	��@�2*�&8-��t'@�@��D�S\�iq��`h{K���f�W&z�O�R��/P��j<W%r(R�.­�
<���0 c9�%Z���^��Ϸ��&�^�T��ˡ�/�ٯ�7�Z���5��󬂃���_ۉ�E�t�o��P�u˪^cq��Uc�㹂�;�{|�p�������sU-ҟ�"�V�xs{-�"W�����IS���T���q�P_6����(1�4�v2>��<�H�&tSὅ���wu�}E�r]$�?硰@�5Ů�A����}}/P�lA�O��G��7|��䳮�#��kx�f�H��%Ȩh������Q���ؓO�7I�fo�A��oΦ��p�o������ �i5��P1*���Z�c��@Y���iqlS;a+=�y�7f[�]A[�sz���(er�Bz.��1���.�a�B���%�?�q��5�R��-��ܜ�&������W6$8�Q�,���sNY���}+����(���e�YVܧ�Iރ���[���^%�4���*�a����K%q�I&�"pg��d�\�ʢO.�C��ݽ(��8�c��HB�����ؽ�r�k��m�������f�(Kk�u��*>W��xYm�O�s��/gb�K�c�q=�;�`���o�$O~�o�J�ϔ������#��p}�CM���q�f/q���_3�"�K���l�v%5�η�r<D{���Ul^0�
�lv=l^�ENy:��z�	���A��Ս��G��{�ɑ���&���ܟ��Ɂ��'������`%��Q�\��w�P?(W]$ҵY�k��w`Q>��!/NS��%8�*��;�㗲J� BO�@DI����h*&3-� �>S�k֮�U)�q��]��;���*�ȹ�?�؞L�iH���IUQ���a0��n��/U�a-Ɋ����l��JS�x�<`AB؜ ��tPM?�AUx9e�<m�Oj��̘��rj%�!q��#���]�u���;�!���HW(��/AB��]=���+(�t�8�i����5�gD_�\ȤW+����ÒTi�R��O���2�kv�=���.��#�n�l%�c78:[uT���yl}�<�-�@%���J�8����-����f=w<�r�QHgq�_<��d(�Y��x���_��z���c�5�Cf,`�:�wI�BT�����p�4ߺBk���e'G"kc���^��q�v��~��sK
G����p�W�(SJ��s��0Gk��7�\_�h���B֙��;a�o��h{K����SA�Lu��$qa��}Ǉ�^��cww��E%}<����g�	#�����_�2��Z^r	*��y�5=��3�(@4�|�b�p��D��=K�;�� �u�m�7���!h?y��
>^�5�r���L�)���a�}�c��Ŋ�%�&��H[�閶��F+���AO�g�w؈N��F��j�2�^L���x���y�����e�ݱ�����U�^5���V|�kn�ǵ����;t��`)U.�Q�Ź$��KN��7!�/P�))3Z���M?�|F6����w�Tk�q�U�5=*�֤yne2�w]/2�kу�)׆�~�ʬ���&ߤAU[���(>j �_�9�B�KNK#�V{-�;
@�~`@�\w�y�_6.=�Z�Ki�:5�h���nmyu�
z��6���/(�ޫ�z�勌�s-����/n!nĨ��N04H&M*��D[_�r�D�\�c&N���d�l��v8�d��H> ���Kp3�?<�K�ض��w���О�Uս��|�xA�n�����o���[��(TK� ��ګX�=j�}��p���o��>BZB�8o�9� ����B�"A�	�M� �Xˆ Y���~,s�:@�ٞl�����Ϸ�����f�T��� m]�ď����%�cw��&\P��JG5�w7������n�:���RZ��]�`!L�~�
����3�|��
1��"^�q�s��O���^!�O8��;5*XLq�����8�_-h 0��?V��Y}03�ʉ��:cV����P��?.�����{4��}�vti�ǹ���$AI���i�"�y<���H�><�d�9�,��P��2��j<FF�Ls��Ntv���Y�Ԅ;3.�\�!V���܂��C�ƛ���6Fh݆*f	J�z^���|U-���Q�d蜑l�(M��7�e^/n*���AG�R7���y��#'	Ԉ1@�,CӁ���KO����k��U�p�?�R��7ջ]�<F�qst��Z�#�X_?DK �o�#V�-�Sl��B

�Rx1[�BSA��|�Q�Z�r�˨�m%Iݰ+=�V����{���<�j[^\�7�c�n\����z;�$fP.�\VXlxVHYEB    fa00    10c0t�.Y��-�D���{�IX��,4���u��}`+��ә�t��	���F�2��|~�Y1�=	ː�Ɲ*��&hH��M�	�8CY�/��CE���ò|���Ĩ�V�xg�.3wQҕ�w�^܏�\�W?B�7�d��f�U�i�ķ-@$[�#���J�\�\��O��� �,]�P�<v��V��C�S}�o#�Ay)��/�h}(�9û퐡�J9C��Ͼ?f��OU"�-����h�j?r-RwMؗ�Ě��Z���n����U�9�f���T��+@���E�\�G;��і�G���d�pdS�8r��"V͠�|NB��FtA��r}�:|-S�O�)�2��+	�V�H$l$�����.�A����Q���Z��}	�6y�G���zH�3ޗ6U���s�wbk�f�(C��P��O�ôE�^n��T��v#��!��n'hV���s���>Q����P�'L.P3��8������Omɮ���q����9W�^X8?\���,�#��(�UJmi<F�`��@��?R�6��c��ʔk������*��}�~�z�5��2��`k��������Ќχ�0@B�쳭�	}F[5uN!��S�޽����4�����)�"3���7j�|�,�0L�ӔK'�Zf��ت�Uuu������$��Qhwʒ�媬~F}{���?@����~e��W��0zX��$�}ϊ�7�a0JK\�/�!ҿ�Y�BOaN2�n*CR��嚾��mW��N[��$��� ���$���2zP�,�Ӏ�Muv_5!�ȷ�/g�v@���qY���OQ|b{���-��?g���l	�;1�u����c;��I����1)�9�kj<�f�Ҟb�M�T����|'AA�$�-n��]B�p�Cf����}�.����H���Y7�}دu��3�U}\�Ѱ��s[2^ֲ�o�^<\ 32����1�<E��p3u�n�U7�>��+`�����h����9]Js�2��,Ū�l�j�/�)�nN9gZ2� �CJ��\d#�&��
�8)F�P����4�0Ek�ӱD�Rᔉ6��g��q ��ۖ��E�q�2��?�m�54����SaV��\a�0֪Ai�}ftx!�f.$|<��6����r`?�U��9v8]Sb$P��٨ɶͶ���9g=�� �(���mn���op4�@��۔Lw�)�E�~f�^�=��<����rʖ��E٭�{���S8(�1��z�J�����YP��O��S��9E����%Da���]��W�U7z�u�����H�,X_�ջD�I�!�DBK�����\i�$�J��f����.oDsY�A�?{�������>�"_Ecg)X���H�ߎ\4�>a� �X�_[�Ñ��}�~s��f:6:�F&�"1]M�f������b;R��6�7d�c�Ev��	
��:���1����rW�[�H9q�Ք�'b�o�2v|QX�����Z^>0X�&�(S�/�H���k�B^�����gf-2b[fm�>��aņ���(�U��JjV@BS�d؎z�G^1T�q��G@`Վlx��cg�º�<�����Ս�^$6��2��[�|�$��\���)��v0&�y��n5v/B����!��:ȍ{Ԥ�I)�e)i���.5���q0	^��>��U{|�[�~�}'��<Z#����N-Jm�h��5�$|VNb<�j�Xm={�׮�!m欂�${G�O�����tD�G�rmqI[��M)@e�v.�)Y\Z!z��Iwy����v�І*��v!��mE�j���{��s�"����/6�`=X	m;G��ga��)\ rG��ĕƱ�A�x�I��D��d&�PǶF)��p�)�%t�z�\�e�0���c�0"Z�/g(�!���4��AHB�M}aP1v�n߯͗��H�<ME��[�z&c�Ɏt+$Y%B�?�:�Os�s&�#	�ߣ*5�>��e�(�����S�b�n�Ԍ�gGB�7�������z�)y�v��	+F/�����&�1<�1�87)�?I���bv~nH��k�Ʞj��&ֱ?L t�!ؽ; �;�<�%OV��=/���{Z�Z�<����J �aaUطH�T�|4��4B�R@{=k�x�������Y�4�L�-�+ȩ��#;dT'v���3(<�FQ3��N��'�`����� 	p��	.T�h�>�f�`/_ϳ݄_G���ޔ�ԥ��bv��!\݊�<��� �s���-�G��_��	�V�~����#1�c#03��搠�Q�	zH��	'��y�V�j�7�#�m�b��+X�+����}~C������x
AY�����,�2�j�;����h��7�W�T�NB>plY�%"�����
��3�&-
"�H��{��j��=�9���	�ܽ5҈�<$��>1(>a�WW�qK��$�Դ��=��\�7N��[��,�i�U"�Qd�i����$��G�gs�o�5-0�7'Bst�BL��惑ƈ��l�An��YoĞ��y5�"޴��I�}^4�&0�\�ץӪ(CՎR��to-Z�X�Y�_ZԒ�A�u�W넧�;xv9	�0���aJ{��J�}u��Jb��b8��q��L���{�����E�"��7B���s��%���=�m��?B=.�Q;Pq֩�O����Y�<4n���d�Ӏfܿ�<��YrTrμ=�Y�Ͻ�S�\���>� etyX-?��64P��$Vj��R&�=���1�-��A��`�gZ��U9#�v��2���#2�����fd�gzP��:K��������>�~{H�%v���B÷l���#6Jg"�rϪ�<-��u���X�H�B��o�.���͖*�(b��O]�w���P�C����p��7N���ӝ���tG��oB�ż�ˠT�:�j���Yʤ�j�Fw)�$�x���O�8��7�x�&�[C��h�pa��'�q`��K��{~o�0�/D��xuK�Y��A��g|���H�N�e�|�Q,���� -�	�#(.�� 0+��X7��8��֋(��c���^,d�*���+银{R�N�{q��K�v�=wq�C��<�}G�R4ۓa��8c�&��&�����h\� ��M:�9r&s/v�oL�qz��v9���|�������(똏���{F�SQ�^�֝7���߁���:�R����jY�NJx]E���Il��J�_X.B�w�x +�9��2��w�L�Z����	}i�*�P�wD�huГ�7�i�v=Z�nK@uj�ґ ���I��"��VB9f���*���oL�Lhv(����@���S����iSJ�̼�����Ai��Ix��iw��g���/Cé�n�FqJ��(<vbw[=�,�ژ혔S�e"��Aױ
omNW�t�F!ɪR����KpZ��+~:�ÿyo��"���M9����i��z� ͯ����7Ӑ������[�tjη��g�HI�>x��tԊ���k����J�!'�+�|`�k�{���i��8��W+���B���ԝ2U?��SPe~�|��=�ƪ�M��			��ұ�ʿ�1�F��L�n�x����/&􄅒1~w,���JO���L�9�`/����6"��ER��L���3K�,�/�+PM��}%��\�� �4�r�O�?��������Z�y�+�����Jo�1�f�X��9%'ۺ�uܤ@�8o����!"hk�仸~[}]�M�[�޵��	��;�O7Ps��� bS?oVV�	�����n�1~��A�I��|���C�r���0we�aCB��粇���_���Ǭ��Vu�"�Jb�'�WSmm_�41�F��t�5��!Yڄ�`�x��{�#�c"���5�f���ݙ<�^�B�2�Ա���%�8�)��B|��ΎLW�01���>_2e�M�ZͰ�;��P��}l`����(,Yg�N
2���8P��'�̔w�23���x�pQ�AKc3�˟��͸F�IR@x[9'P,B��hh��s4�+����]%3�E s����i���� tb��C�᩵���-4y��sX�:N.��L�[o�j��?	��#�o���'�5hφ�Q5-Du�S������C������J�(�2@���@AC���[~~�Xs�n=·�D�a_{��şGw "#��>n���A�oZK:XlxVHYEB    fa00    1140���@�ɖ�M���١���XZ@j�ۧͶL��'��qAꑛk&.5�������*|�uh>Ь��lU����5���8��p ��͘Ph�H�{E$�����T0�z'M��hU�A�S��㚘��H\�y�e:E~8yv=YGo�q�`�C�?�����Knt8���z/�<]�8^�k9m2=�3e�1udC�s�UC�7�
�8n1� u�>�h����hH�J�6�W��n��ˠMl�Y����c����A}GI=�kw�xKf����H~k��Y�Ȱ!H���=�UH"w��/�@*h�Rd�W���,������(9�"�Q���" v��*q�`M���I{��"���;i"�h�����\]�l���D��"Ò��'?]�Ln�����~x����$��X鸞h/LB�)SC2��57I���oF<d�T��e��U6U�T&)� 'R,�{E�︠��⒔Q��WQG�	��~��֭�SA��=F���(�����Fʃ��0̈ۚ��V�������󇻓s@n���"#*E4�L�-��$���%�	�Zd��Ss�駯j*wl�׃��>
�����+ �yò�\��_��%8���!P5쉟-d�,�/T{���t����1Q\fiG#L�g����6�w�U(�Nlr^/f �a%/�1M`4G܌��ѫG�r�Q��I*zoȗ����+Q�Nd�i�.{<�������̴�N�C��⭒���Ee۶����<���LՒZ��A���h^��LV��rݴ%7
3؄L��ڵ�P�����q�.�xp������7J��DOM��S�MqY��ۗ����9��[L�
����
f>����t��d�
�jM���0dP���L}I���ӖsDK���z��Xג� &J�I��2�J����;S_�lUZDVV��F_B6�o�a@a/9Q��.[1Uxg��r�"^t�S�'E���.VZ�Vĵ�G9��.O5y�bD�,�=e|Ed'�hS�����r������&j�KQ�9:*w��rh�kM�5�ub��Ӽ�5#'�ž����s*��PĴ�?��7�}0'�e����&Cm�dQ�cyO\��(1���H�a'2z<�T��k#b�Ԋ(����D*�:U���|d;u]���d}�E���SǠc�o)�;�sy@�r�QH�����J��4vwS�VN��H[���P���`�>>:!L�|��K;0�C߬��ǚs��w����������C�Dl�%~Y�@G��k[���7�/U������!x�[��#!�	�@����U���F�"'d�9u�RVEK�\�"�Vn�0�/��+Ct�]g�:4� 
���;���id���1r�.0|���#'�ѝ/*F{�yJ�th�W�s�Hu��<Y�����X�H�o&�^4��<z~���|�&,��b`�O�Osᘷ���_�4m�Ŧk�)\i4�$�l+�녤��r�9�D��uӛ� G��% ��+|l���Y�A��	�4��ua�_7����a����s�H�=����Y��Tj�$�"Z�C���" ����r���P����*y��[�}\1	�Y�X
hj�V�3��ex�R���sx�@G�1fLڲ+�o�Ն"H�f����f��tWOc�NP_���~�>��>�n-\LeF3B���L]p��P�Q\�,A�@��bDU9a�v��S��|q�ھ�ڿ�I�CE�Q���Dt�[7к��(�`��:� 
 ���ݏ��1`{�J����h?�	��ʝ����9�}\����o0�M��>�?X ���9�z�VI��j\���*�<�4�j�)9j:��a?���z-�J�u����O��7WH�(��ӢTee݊T��3��Ɨ3�hW��n���U�{����\�H.�C�귷I�W�$!��O�f�4+���zo�ob$��n;���BK=Fn�jp���O�qj�gp������ԝ�ᰍ<���h��u����%P@H���U+���vf��fR!`7Rw t��^��4��c����"U+�H?���.�W:P�1c�H��Lҏ��̂���Qˍ�V��=#�Aa}ҷvgZO�%����Z�.`�-��x'Xc�p�@�W#P�����<�����;��������H�E<D�H�Gud�'��f�	����&�QUWeƂ���a˯*��+R���u������:o�K ̊��B�I����22����L�L�¿�8������{w�	
��>���R!���-*f.N�^�v��ϣΑD4�2�] ǎs;�
8g������8��G@�'x5&��$z�*���dI��v[���<�q8�ft��٘���!�P?�X��z!��2�-n#��4�}TÝ�	��n�钵Z��� Ա�Z�O]}̵F��*M��QW��ǁ�t��*���A�����Չ_�� z�o��V*�/��y�p����~�B �9{�M���@��F�;��9P��Rp���2��p��!�j���!�& ����w:J-k/`�{hƶ��V��E�dp<3`�����4��q���:T�p$,��D�摹�֘��G�\C��n�M^���3��$�X��2���Zq�.c�x<�7�U���z3��{5\5r�OX�`h*��֡Y~��	�U�xmz���S2��vǸ.��+���2�����F��C�����Ueo���������=�{��b�9qI�	nIQ��Y�x~����E)��ӊ݀Ņ��%(�K��e�JI!�A��!ݜ!!&����}��6�k�2�sp]�|׃{��+E���8HӞj�P���Uҫ�����i�����N��>Db��{i�s�M�o�N�lDh�OS��D�NP��r�,C�;����8����2���!C��3i���6kw�S򗷇t�'l�{��V����qgͶ�j���K���N
i���v���Mȯf���ؤ�.�a�0�p�������ꩿ�e���l, }��ܚ+�+<Y�|��p
�s�� 2+��s�OE�C�{kܐ�
�[9·߾U��>E2˼��":�A��YBk tUǻJ���s�m#5�]8}��P�*����0 ;$�E�_�~O.�O2E�u�Ö́���`6�,p3�	Lt�o���uT�4��1W&�U���zl��v�����B�+�Jpib>�7+g׿%��r�����R��v�k��Ԇ��Պ�t�o�mlS��� �B�۵�v�k��0�Y�퉊� ����}ղ7�? �>���� C�#�Z�iF`�)�:_-8�op��a59����z��`0������"g��
�(0��
)D@�N+W#�]�7D��0�<�>�v��=n (���Ǐ��_Y�^1����a����Z���JW�£���6����M��������&i�_eo��cM\�;eC��$~	Z�閜P�-���wM6����Pƈ)��h���~�+k�F���]���K^Y���$�8t������p@2H��ի��p����#JYVϳJ@�:"��M�
�K \7_0�e\N:O�,.�g�at�^;��WB7������c��+��Mk�I>�,9�J��Ҩ�t@��Kq�t���^Y�a����B"�/?��W���՜<��?�ʚ�و�[ ڕ\�zLi� č����j�/8�6-WC}3��2��x0F�?΃�Ȕ�D��EC�K�3�У������N@[�c	噞�b0T�[6���?;���Sg��M��N��\,A��	�G#"�O�9�:G�����,���g~S�\:[2F�ɕ�x�J{C��$�"�4o�N��`��d�^{p������Z�l>o���k�t/��^��/���-B����ð�-qę�c�P�a�_J]7�~�h4�S�Fٝ�������D�0��S�AA=�-7�� Y@��]��d�`�\�p�&�z����q����F6W7۪ӄP	�g{��N��|�{��C��gb���7�u�;1ɋ��t�V4����>��qvwW%����X/~�6�$do����s�3�{:N���Z��t<�^�8)o�`s|"i�\�iܰ��<ӂ�l|��X���x�f�/�u��r��]�S��T�y5K���#�ȁУ�3�"���=mAu��կ7-�XT3	�Rb�z��J!�z(!g�q#eIS�z*;�|���������".!���^��0֣ (���Z����xl�P���S�!��P_��mt��*)�� }��ȆŰ?�!��@�3. �a�J�&>��CU95(�TMC#5�A~|�P:��M>ǅpB#F��L��GCe���U�����\��:�0_����4A���xmF���l��%��C
Bk��=XlxVHYEB    fa00    12e0��㔱��6�So ��ǲ����ȓ���ܕH���f�����h�/�{c �ⰶ
�	�mД�-�B2X��֭�6��)�XJ=A���DazK��[�D(+s*�}g�4�6n�艓�AT���`��;c�/�i�(=]�y��?�'��-�&$@ؼ��n[�tLeN+�[��R��v��F�ʳ�c�<�����a�l�Ԃ���aY;�"'��P]��	[�c�g]�jM7�I����\�г��O�-�է����h`9���+���7�.��z��nxC&"�X3�O2HΙ�uaOFX�x�f���A��T�26ĊHD���xf�)�]x3���V�����plP6��'b����w1�^�y��@��h�B@�K��L�2�����π�ʘ?�G������7-�%N��D ��z�\I��n_	��U�l�O����ϖq�ƞ�^G��KX@R�^`{mA��N�pg3���{�ڵ�I����&�u���&3�s>x��揞@E�eb�I��%�ڲ�7�,�[i*g[6=��?6e�А�JX]�[D1ӻ@���,�Oԃޛ[~j5DM����|��O���$N�r��P5V�E�$�q�Fc���7����f9F)����f�v��%/�ؓ����j��q�k�m����}dÑ#�[L`z!�*̉��60G)�1��;Q�$����3v�t�@ȑӲ!�7b.L�i'&�/c���
�9�=,��NM �=�x�~��G�7�*"aF2��9Dz�Pbv��;�ҪH`����gz�b��H[��e5��0�����P�T���SF�g��*��ATӲ�����?XԺ .����q�M���)�&��]3ʵ����9�F�C�ɬp���	�ݛ]
g�"X��(���=���rr�=Ɏ!���{3P�Y�L�c7�(�(�&��h��g�S�lB?���@���{������hX:F�Zm���}�I�꽩ga���2�C7�����%u^j*W-�mM|���M�!e����={\*tޔ�d��/jC�ˇr�w��gˎ�S���a��"���}5�1:��ʲ5̫�E���0���M��+J�VU*���O?�}+?��t3���/� K�� �aP�N�"M��|��ܘ�BOȔ+�7+��E�~dN��(� V�"�W9�;���</Z�Ru�j#�rg��7c63:ikyZ�#��g��XC�Ko*���]Q��� L�2s�>e{�M������B���E�ߚ|Y�q^��>Jh�5�
c)�����Dr���A����|��u�k��;��|� ���2�f�[�Q9�0sR@�y��T.�:��5�5٫	E�*ych�|�I]�:�AB�'j�L��Ou1T 	���V�y�����e��Cē(�!�}�S�I�i�I��d��J�UE�J#�ᝣ�G��.�LU9�����PL�zCy]K��S?:w�꽟���������#CA=.��R>I���J&LNzR��W�^@�u�Z�A]�b5��U���������i�0r���?Ԡ�PU�j����
�
������Jg
g�P=�XnK��͘�  hv>!;�y�ӏ��"�ʲM�����N��s�����s���I�˪���,'b��TQP�l=tE�$��H~a �l�H'�d��|/ �d8V<�b�6�j�T:�),��5u�:�/��Kê��U^��6.4a� �zR�����EyGOj��r"}�
^z����R-�2�$ 8#x�F�Qz�<+����lt�"V�Ì�R�Ng�q�����$�g��߉.t���3M$�5kD���y�X�À+�LW�ĔL2�<e�<(w/��g|�	 {��W�g4o<�Ly�O������a鑠�	:B��i2�Y��
<nu>	�3hPKS��QQ
��E;)�V�[�t�2�Km��u׏�l{���P���λK��C?���?Q���A�u���b��$LA�=�GX��4�k�D5��G?����0�j���8�:4"	��$��#/)t�g��W�������m���i�0ɣ��@ ~�xq���|+tƋ��w3��j����e�F�T�)��g���x5�zB�	�c�6��y-�N��o~�T��W�=e����b���-�}�{�T?=�Z_O���i����YY��tk�i��#f>�AU���넑U���X�`ɼ��x�5�� p$�D����-&�lȧm�??3�*(h��݄�#�A`zZ)�����j�	0}y�B#�Uu�5O�kZQ J��h�����V�h�n)�!jT��$��g5ϰ]�D��*���K��ϱF�n� ���U%r��T��5���-mȫ
s��-�S6��t�=hl��p 1�Aቻz9��|љ.[��0�kب��ٖg�5{J�'�$�G�l%��8s�t��5��GH����Wmj����ڲ���0��R�X�] K����{���M�9�VB��Ӓ�N�jZ�0����I�,������\�A�c�*��3p}��#IG�^��EoO� ٿT��0����q�9S�k�����4��Fz� �܃F�V�� �YS�;h���2�����Ie���v"/c�g��"?�
�5!?@
��68�8����u��hs��)F��� 3�蟨%[6�8�D���r��r�W�%�׵a�*w�B�=���8Ͷ����U
���}��v�x�Jؒt ]�=
K����\Fv�?/��L����ˡ���/�%�AW�wV�z����P�K���9��T_*�짪���?*�8R����.��7P5iQlBm3z��;]�ۙ�`���ʾz澴���N�����mSa� ��P��F��#�G�w�Vu��`�f�~��i�zTh����@�w�=���D>\�ݎ���ܔ�):����]��Iy��erqN�u�ܶ�Ʉ`�ER9txTp�#/*2ьy7W��yIu��s��r�m1M��T}�W��_��~V��������:Cp�摭Y�͉�j�<R� ��g{>w=�[ں��7Lk�`�w>Z����v �0>�&��ס$q���;S��"Y�/���L!a۹�8e�/C��c�Ӈ�����3A�u����;x��r�d����>F����-�$�D �=d\;�91V��θ�H�D�y� /��b��pY�zdt��- Gh�Y�a�p�
�������R����J[Xq9����{���H�cpэ���:I	�a<h-��AzD��'<iX�ٿR��^T2�7!���>�^A�/"1��@�����������z��S5DL��r��E���]�ʒ�xEo�!�fQcN�pH��)��fB�Ǘ����Gi���v^��Z�/�X��%}�=��nj���zJ�\�r��nt��;�a��xy:����(&GQߺos����m&��񬉔��&u���"�;x5o:�
�ɝu�]�*9
s[kV6?o����*���v�������%����^�ɮ����-6��*�8����[5��A}M�RMx�s\s� @�x�p�]�WH�|��X�q6,���ݨ0~�Ĥ�$��^�C�n��Ƽ|�X�Ne4�U���TF�U��a��Sy�:R�3��?nG�:����Yը���R2{�&��3-������j�H��(�:��0_�{f�ܞ����۟$�ַ*}$a��@'�5�I�t�F�SB6��<���G5�sKnYYƸ�k+9K�CMu*��T�~��]^CA�R?jf{��Z�p�ao�O'���f���fN�g�s"o�:7	g��x�������D8ka���Gd�5@ʤ
���46�٠����ݐЮBQA�[!C��/Wh}	��X��+u��"s�nŐ���oxK�}e� U�	7�V���nnp�B4�5{��w��@��Aʗh�#��'G�m��h���"�UPp� �� ��8�y��v�t����\}%Ԩ0�艑T���ߪ�$
E��C]� b��:t�oM�u���c���B�C�J��"�eq�)w��#\\�1���o�-�ከ��X,��bc�0]\-ʠH����5��/k��	e�	���[���
V������z��_i�u�C�DbJ���2Qa�T5���7����'�e𵐥�벟��mod,ë�Bs:���Kd/�h�:�n�:�B���6���@S���M2±�5��E@���+P�����+��
���)t�H�!��oE�#n� PZ�r�p�M]�Ep��_dzB\XA�H-�ǞD?u�ȴ�Zg�g�~G+�[�%�������`+��z�����P!'�@W��ܜ�!6�gX9��L���笜���$����{�2��4�qE�y�.UBG�ԟD�� b�����;C[ ;��.q�)B�H4ex F�^��p	�\�Z��	Ҩ�:����^�����JG���:��Ϛ3����Ǉ��b�9�Ն�S�R�`�,Ko�
�,���I��>�K�	w�s\i��?9
0�@�\���|�bLd���� Nde
%����hg�6q�����-��cZ]�EA����4+�?��Y�-���S�$]��"M��&�y�F�����)d܊(��&�4!Wʧ��W#����k	P�mi���^,=����'@<#s���Hf�
t
ˈLk�@���vT/:����}?�<�o�wQ��ӧĞ�L�;G;�3��a��s{Z���/���t��7~}2�R�9�n��+� ��P
4��XlxVHYEB    fa00     f50��f��⾚[�-}�Ǫ��n�������en��S���"96�uU_
`=b���|Ojd�K ���j` W����=�B_�,6E.�(nub�6��i�,���>$�ĺXo�4�e�*�D������(r���,�T��I�TC��5�)."Y>�`��/�S��D���Ȣ����k�y��>�is|�&�-�3�cN(�?��8�i�)3l��S(�c��*�m�ef谨V�R� ��wG�����bCT��[rq����H�kubb����H�G�O����Dp���������5�W�D$���xkֆ[aD����D=B��uԷr�n�ą��U#q_��p�%�!�O%Ӥ��Q�r��+��p ѻ�C���-�I�D��~ �:�0� ��?r�I�8��9�<4���uk�+Rm���"}�Kl�j���r���̗����dǡl@v��Z8D)pr��2VSp=���d���{M1���{��t���8����ZGY� ���{Vh��_����I�r�+}��.�뽡��wY�_�x_ ��A����6�}-�_x��|��5[����X=Eu{7s���&���qY-��ږ���g��\�o�P	��Gh�ȺZ�������s3� BO�	�J�8��h=���T���(-�Wa�U��.V���T�-#b8��M� �GQt��� �5(�g��yǷ��B߭���X� �
6�N�'1w���i5��~��j_��8�℻Rb��Fh�C1`�¼��W!�DU������4 �����b	ma���t�4�x���r�:�Htx%d �=\Ɔ
͟Goމ�%,zҵ(A=��U�8��EɌ�s۶<���=N+����}��\r_����i6���sz�!��VMfma����2�]�IØcW5WV<'b�<ܸ��5���aׁ�"芄���K �պS�l���yA����<B�^Lאp-g����7��W��M�%�zw�v!�k��F������	KM=e��!�9��,�X��y�A�(ej��gㇰ	��w*�s����Y�#��8'�kg��ˤ��:��ҟy�M���l~��ؑ�~�'n�3қA�̬5�������k�����'�k}2���.6�BK<'M�hnŉ.9�ё���W�?���C�^�̔T =Q$ۧ8��8=��2dEȓ�(��B9/#�U���kȏz�K`����7�J�2��)AjÒڒ��j4c71Z�X7Ie�[#N��2�9�"�峓���ϕň���<�zP ���K�5u$��b�B���A�)%�vf�EM͹�>��P�h�����xP8���o$u���L˭��Mtu��rßL^���%+�կ�b����_ď��+���������5h!��d޼�'�1!ص�ټ���`��so�3����'��Br8ؐ�S�� <�D����6��Ѵ��߻��������_Wd�Wh��^�~���A��a��b$��ܤ��.kS5���X�2��/ϸJY�<��8�(h������BlZ�Y�mp�v�����ز��-G��=C}���"qq��+��e���ȼT�8�_FYKk*�Z]z�3�u�T�@�x��3�(�����h��j�K���?�Y��\�շ����Rk�g�(ӟ�E���ԖM0\z����;��&L
����`A��aw*�B�K����H�̃$�o��X\� 7���J��:�b^b1M�ҥh��T�<�]�\i�q6h�������FPN�1�μ`o�����]�V!�������3��U0��\����D�/�/J�"��H
���1�ZTt�GV�WN��
i����Qas�	 i*�3��r7�����H a�A�DB����5'�g��? i��
ȑ�V^��>I�'[Ih�еƁ��e9�Ft�0ML�2�� W�E���r��\����Jc+-7�Y���:{Bh�F����NE��ڈЙ+3)����w�2Y�&��_����_퓧f��"!k�!�Q�P�c��İ�!�)|)�T2E�\S��Wbn
��,L��xB��<p-�<Vv�%ǆ ��\�[ћ�u������U�t$�/����Z\t�]��ߢ�?
��v��	c�!�ڽs��,"r��zm��$1��!�P6�y���+��yc��EB*!rք��'k'|��Z?S�<��Y)�}}'�����&��+�
�j(�a��F�,��î/�э��Q{Hp��f�9��}jd�5�VjG#����ϾF~�I�y��!q�#�����v+d ��/��W;�&�����I�Gv��"֝��>���W|��/"H�Оa��t<3|TZ@���:�!�^��I|�ľrrn�J��4�yn��amn1Sew�]T��}�6f�>Һ�혉W�;�Ql�ࣗ�oYK��N.shʹ�U�<Fܚ��N����f���S�of�G6�O�� ��􍗔14�n��_�.g.����7�Y8k�Unn�h|w­�(7��u�1����xB=�v�_(톻����yH��'�R�	�����e�0�R��A�	���F@�W~�Q���9����D�����a,�_�_i�l���p@�~�)�`�VB"���d���FӇ�*�*�`7$5�`�x̂�JM�A,��O�Q�g@���	]��UK�o�GIKM�1�m�鮓�{���^��1Ȧ�|���G(�:��vo�V��Bё?-�"���~�b�Ű�S�>k�x�q�0ݑ�ǖ�	&��ʔײ%���-۳ÆjT}<Rj�(�s	���b�/9mv٧1|n�q4�E��\);sC5E�|s��B��7>���SH��=_�m��U�~����<,���X�R NP��?ҿ���[��M���%�&;o�1�/w�J�ө+�k�3�/�0�6sH�*9�MK�1��{��T��kd"����?�Պ_��hp����*ŶY�HuⰯ���H�'����{�r��Wv�c�&��+�zYWȃegq�)��1()�����?8 ��|��7�(Lf�7y4��x����q���0��-�7z)�F/ �}m��&n-�5�4DA�u��#�p�.����d>�׷`���<���y��͕=�ԽtNOL��(�����Bݙڜ�����D���5)��_�w�⪦-�/I��,�%�G����?	�T� ���&���u��V����<������>|F39ꓡ�1�QR�5��j�T�d!AB�kq`SJ����dT~�<��5��w/fnc�dL��4��Z��a���[I6�'=B����jyy!n(�>�nM������'Y�=����L�Bgobo�B8t�L: �����Z��7� ��K��^�?�b�Θ��9��)�����h��_�\ 4�t��J޺s��S�4��Mi�Hf�N��/�E�V(�t�EQ �D`ê
o�d��o��O&v?��F(>Aԛ��J��6c�ϐ�Q����z�Ԧ*��2d�+G����A��5 ��,�q23d��4�j�Q�|c,~q�G�/���q��T�6%D�Πlq���w��sX�;#ȗ9]�p�oR��@o�W"��C�0Y�CF��"yc���F�0���6�+E�2z��,m@�9��.�I}�@]����!!�I��o]�&X�7����ä����2~�>�F}�&[� �\�Q�p�����7+�沑��vDVꛤj>�=�Ǖ���c��k�@��I&fc�+�y�B������pU[*CM�'�z��'���ɻXlc�+����b�@4��z�>.����u��MD\p��=e,�!*e&m��h�,�b��<�xa*�
�IגnWE�蓵\�C����<2t�)�֝t��XlxVHYEB    7273     5608��хE�3U8jUj H�-?��B#���į�a�S`y!Cq�iCzE��=�d��Ҳvr��sH�a�H���.�`c�ax�:j_�9���^	�p٪�c��Q��8��LG�^}G"ry��Μpg�w�Z#��r���o�z���ab�|�X1�n�Z�e������TX�+�=$^Vt��'�c���n�;�7���Oޚ\�Я��eH����ݙ�^�h&	��ax�jzv��z�a�+K�k����u�������{}#p>>���B2��l��јL�6�4E��
��Y��
�K����M&�rA�y?Q��W�ݨ�$S�R��`؉��X����2q �X��f�mͩMo����R\�_�^f+�:i�	cu�V��d���wy�w��I���ZN��Ғmi(R]g�d��M��ۖ���e������
znJ�}�^��QC�DQ�7� IL���h�KO	�;�%�5���&��˶����x��]qG�� �ǒSi��$��p�h
4�˱b�ʰbcn(��:C��K�$ d��([ѝM3[3�dҸ��w���K{Lg�G�v�	��rq8�q�H��GvԄL�p8=K�b6����f�iW^T��]{WS��z�C��,��{�|r(]V�K^6��T�����F��P�f�\~y@j�4�(��V���[�5�@�~>xT�b�2���j�~�f5�q�K�z�|uV#V[�(�o��0��R,�#�N�!����cvǒ��x{E�1�1L|_��k}��Ml(s(����L?V ��B���U�ƥՒ("��k�b}|�}a����%�m�o��eӖ�b��P�FNya+T�{�٬�n?D5��dF#�*�*m����5�;n:�K����u*��Fa���U�^H$�Rw���B� �5G��� N�G��������Xf�v���[�{���i���Ӏ(LNT�N�:�Eρ�@�����t���e�y*vX���Y?Dc`��>-�����i���?Q1�´wgU�A�1����������,U��.T����P��~�.�4���eϣrG�֯��Sj�ƺ����P�D�2=2�A�������B�ʔ0e�����]�~�����bg����m��(�uꞵ�qml�f���H�G���g�C��ԧ���`�j�P=��/R�Tn�`t��P�ھx�Ʋ�^18�Y����6��Ԝ��_�{��R�(bzM��^:f����rs��=֭O_�D��/��{�bG�`Ɋ[��b��*� ��a�$�wW@Tr[q��uj�%���Bj�ü����CɎ��4/���p��D�٘F�&��|�]�'!�6�