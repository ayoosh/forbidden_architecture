XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���&��l�) jV/�O�G%�Nha� ����b4A��2��(��Չh5�i�C�I>Ŏ�I�웶��n����Z�$ ��a�L�;8~�B��aʚ�\�_UN�3܎O�̩I���y����,)@���`d�	�]�OHm�7�is=���b���Y�_7l�FE���j��4��n5?$��P�*���+q]�𯜜ab"����;ɿ����%u��߷���SÒ��)�P(I��K�o��2>�P]{�|}C�c���:��?�Ď V7�m�²�������θ�B�K���o4���f3��(�/����!=;���=�6��9�Fk[���sr[�����.	�z�
(�7�y��W���1T�D��{��B"���8�m���݀�6%�KR���Mb8cq��-
(�F���pm�A��h�$ao�v?�~2H("(or�Nm
h@�C��ۊ*���X������j0�G!���X�:��"�>�v~`dI�U_���\�1��|����Kڙ�nE!���K��Z<�}F
��x|SD~2i��;����cy�G����~��t�X��A7A�lX\y�lJ�zC��o���<�6���p��D=�2�����ے[�D�χ��3~J����VY������:n�q^ndU���=vxݒ��CL�hq8K���b�����ZQl䢧[��n4E��e1�PWl��ҽ���V۴3Sz<m�d"��uIܷ�ۊA�e� �w���N3�hڶT;frXlxVHYEB    aa31    1e40��w��h���2�R�,�E�L��RSD �z`����ŢLv���"b̔qrc��u*~Z'�k�~��s��h���sn�|�ӛQ�W�E ��n�C�s.�(�xfA�������Cs����ķ��A�97M�8��������_���^���YZ�R��()j7�(�O���+���'ȃ���RF�1f��^����;Q ��GT���9��:ş�aس��y��`Of��3(}�2
[U�0V�X�U��wS�o����N�gnsR��a���?YʒQ`n�Fק-��?d��jjڄ�^19�E�8}[L���K�.���ގ�!��`#�[ ?^(�s)���[�ed�Vd?�6{�@ �?I6P�[��`9����wםƍ����/ �f�
�J�L��5q�2Z���n4��iH',@3��pKA�nS@�ֽa�K_|�63�AmX�b�$c�ۛ�\��5��e�ǹ��>��'p9��M��Q�E�b�~R1�":�Ml���n��.�@���sEZ=T�%25��+oAn���=�;�^�@ �"8c����(���q�k�	_�	����ԁ���xݩʽ�{�+> Uev��q�^��*�:�~��R�q#O��L�! 9����/��S���[�2R6X,�'���3�Us���v�m�$�N����R�c�[����#��8w21�9�DS�.�ԞgQ%ܢ��i�wHX$�҈��ϸ����W�`����m�+�p���9�eԿSTsq��,��O����M\�*�@�W=���ߊ��l�R�*�k�mS<*�y��N�OP�sX�t��DX㖢�����azܬjq�ˡ~4�.c#�����6�[?"�(���r���ҧ3�{��ؤ��T��zNV�qL��mKQ�ψ�e�%|J������jdh�W�3b�h5��a���&�20�;"����ZvD+�J-��	�ЀL���Q!ӥ}������1�m>w/8���x[�ov���bͬ'
;U��sE 5֌�I� �l��7�67�e���)6��9��=k�i��ˈ�ƀ.��a��V�ᅪ��*��8,�,�����B!xc�l��*��%�䣭/�����Q9�bb����Qj�roE�H(јt�T�H�dY>o�4R���	�����7����6����8�&|�����+���>q�t��ӵϸ6�$�3��o �J97ד�	s>5D�B���q���N������,\�H��/���5U���� `Iv�4�O_���tD���}�K?�������Mͫ�N�g���8JT�Z�FW��V!�)���o�*Un�Ċ�Vhg��*�e󬌹����6N*K�K��UA������y�viS�;{��DnsTX�e�2>f'�R���b��6g�mк�G�b�_P�y��c߈�y_,T$�@`�lx1I��Q$�4�*��g@��E�����4�:>��6�S�
�a�ޫ�=��I���v��a�{�ϼSp�u�O���S�YX��l�mYȟg��#�^G
��0`^�P�(nq���Yz�S^�
�B�(�n�SɊYm�V��߯b�d�iMR����qԴ�hV�*Ɯ���O�\��hV'�Z��(a�h�~���@����Z"��/�!s��HeXn��,е	����Ƙ"�lJ�Sx�*�_=��]U�|�6��ʹ��������b����)�S�&۪�
�*_A�;J�����6��*��
s+@�[)�h‼E[oZ���N2���R� � �s��Jzt420t �#躪b懊�L���0��1)q]�;��2M�[�(^5w��\�·�(�.2Jvr ����[�(�g��9��I=3	�g
�pSc��SR�eDB�\�e�z��+�u�f��u������:�.�"p�&�,��W��P��v1���<���6+�Yͻ)�է)�j�,)TRS$yѥ"�wH
ʑ�$��V<�����ۯ�X��k�6~�xDqZI\Y�PD�Ɨ�����S�����nkt�&:N�'�G ��S�o��	�-���s|aĵ��0���ʩ��f<��U�����}� ߖ��~�_U�l_���Q pMc���锃�����X�'���LK���G�˱�R�9f��F[�����
ѩR�>�S��)�QWh�A�<o9k����Egl�i�sWr��6�z�4v�a�E8\�����O%�#å�u|ن4���:-��¯����0�w�����/��}@�J��\%���@a�rǁ=8���V2F;��0�x���]S��`YY��F���1�:jssw:q/�q�V�̰�pm�q��6ja_�;�4�����C����չ�/]u$_�ϯ��RoB�ƾZMo��Qn���ѥ�AG��Ո���ڬȌdxZt]��±|q̔�s�uߖ{̎���DŞc|��e����:��Ϝ�R*��+<���s��^盾q�[�l΅f޼3B��h"���;UI�6��$���~QT�A��J	�J'�h:|�D�R�Zk�.F!�?��+�V���iW��k�f3�"��>�NS~t^��Ǜ2j�?<lŀp�ð�U>J�H1�rĿM�I���B:��3�I��5g��&݆�hǻ~Aj���)K�� ����#!��_�8d`-���z0W0��5�x N��C�ԩe�8��?(ʬ|��t)��\xFש*8Eu�m=K���6���1�dh�$f�d�S�޳̥д�vRɤ�?� ��-�-��IλW/��p��)i<�� ����?eVf9��UV�n��h4���4oKC3��m3:>Tه����Ğ��]�{��N�L'9���(����B�����iO�%�D�n���cG,�kR�"��F��Z �/�ǿ9LU�:R~�K!��~j2��my.�}�kۀףm��6���vJ��p6y�+-�hg��-�{��i��q�+��(
҇��}z̔��Lc$�H3;����CX0�ۅez"���I,�N��?����oe���y��\�OT%�K\邏w��j�>w�蠆�E�k9F�43 ��qW|+zM1�����1D����ZY���Kǂ�kT?��ճo����Iۄ�$��%�i�Q1ڊu���5ȴr�0l2��7��x���]���%����g�X�\�i��]�Pd9��=AZU��n��P�n�#E
��e$K�_��w��b-�����w��{�9�P�������/�u���|�Gz^�F�k�/;M�kQ���J'jS����NX��V��	��M�R6�爹��(������V~@g�
R�����-�ѱq{ʍ�F%��p	�ۆ��AӆJ��G�U�������V�Y��϶͙��4�Q�vꘖ0��#T�&eQ�3�o�:�6:G�m8]�@��"�t?�}���GU����3�eZ߫z�#�D3ƈ<�n}��0lub��c��q�p��#F|Vn�N�
%��OaK�G�K���-��W,�2���R��P�S��Fϛ�xT`Ŵ�)��k �KĖA;�H��+y��N$�%p�,���c`�a&�Zu�_6W�,��g�J3�b�N��Ydt���	��S��-���K�C^A����K��6ÍGE(���K-�C5 ��Ww��U-�?�ڡ�r����o&`k>xٰk������Zc�Nn��|��� q���ZKc�fB��nMG����`(���5^�����3��#2�1OIX[X.��]w"%�fa-�{�����L4�n�P5nq.1����Y����e0d:u�ԑ���䠒J��/y�� �r;$P�Q���忀����VZ+-���IM'�Bt>�� ֣���L����Ya]]L�-����`���ym��3��K��8^]��.�a��Ov�W���M��Z���
�25Ӂ7S�-1�+�LЫ���/������R���@��w���R{Z}Q6D��3���Eȟ� ������N;`�I ?˰�yr�
�.4�؅�ej�j�)+/�^�ڱ���b�^���ĳC���8�,�\E|E^ ���]��ת s����4��y�9��a^�Vr7\�ǏY�g3��֦B��� -���7>��9��h�Zo��ʨj��M]�2E��{��:S=-v\���(�0"��7��;S�γV�����J�	�M���g�-(�[L�T72� 2ސG�7��]M��"�i.��H�S*	����Y(|�/�]SK�~߇���+]��v�)�W����VoV�0kD�,��*Ӡ���皿�be-{�Z!�I���?ml8���!Z�ӄ0,
��e��Oq��G ��n��8~�����kk_���]�-�Л�.�@Fp�1�9e�I��g}�۰����;��1	F�5�-'�7�2#��&�>�m���z����%5���6���Q(
OP̶���(C�_�٣�D�@�?�oE:v[�Z�n�Hf�9�*r���B�� 0�8���l{l&�����+�@�S3lkU�`
l*o;��<�ǭ�$�s�}��&��mQ�<p���|tD�����#=@� ��@�_"�0Ԯ�fl�m����[�V<�����|�/����	�NC] w��3ʂETM�¤��p�G5�����_���&�7�}?�Gɔ��h��҅wC�/���%���1Y�I�p���j���
���?������<�TC�Vˍ��\�\�(�UD ���S���J F�1�� K�����7�SOx��M�~�j�(
t�~���G�����2w�}�X
8����0`˰�c��#��ʮ�|<�v���3�橞�@@���S��yV;��Q0�=�ގ�|�B${�e�l���e=i2�`16B�[�{�	 ~t\	�uu[��&tm77��ʎЦ�'xk�5Uf�����c�Z	��f�6w7џi2H�9����n��%7��{$��wSN��'� .԰��f/��~?Ų�Tڳ+�,��wnd$ؓ(�)d��"=��o�eW@A��)ί	Nh�������k.�R_B�h�w�l��G5�*8�zy�jiG�|N(��%`�(R�?	E�{�?o��x%�~Me�x�gtE����y��"�c���h�6����?R�=L�y��`ZL�q��h��:�WȎt��)&5�~����$�'�z�-�JY��Ke���u����#� R��JȄ&�a7�4: (��qu��Pw�����Z��e_��!v͛V���5�p8.K'��nR	�����0�����*�[4u��&R+p���w��_��H`,6Fu �&����n�������W)���������v?���2�}�Ы�U,�|��1�H˓��Ks ��͂�m��қ�C�{���Oլ�+�(��?K�����u�3�e���Q�aE��Ð62���o���; �4��%�z��(���"�Ш<'/��<�� �����W���ٱ7���/k��8	k�^W����&�XX��_��g�)CӃq�� x%�D��@��\@+�#��fX�Ƌ���h�%����+���rS��P���4@AV���Ig���V���<�2f���FY~����PB&� 
<��Y&W��)r��2:�BP��X��{O%V�d�V���"��ᷦ��2!~V�{��Ѕ`��$t�ݥ"�r�mռqJ��n���w�;'����*�|�-n�<�F� ;�-�ȕ�i�T�����[o\4�p6ߘ�����<?w$�5:�ȝ�&�h,���9�*�`�Jn�g6��w$�"���г����P���R~t^��N`�BG�X��`�MYTŶd��>���FB������;z��l�H#3X�^7G���}�.~��[���A$�O��YjII��^􏷛�k��\ē�N%Ħ�;��RO+"���@ߔ8V�š�w�}p��[�]�L�]p�fb�g\��C�[MF�.��3���J��Þ[����ԌZu�o'���v��	��//�;y���7�m�="��$��#��X�����	rm��=��.�wyxQWYs!���u1@�'���)��,�}8R4|w|2V�
�$�<��8���RQ��I�d�۵������$�0�K$�؁�\�!��ӷ�wl���b�����w��&��j2��o�S`,�:��?5��>J��=�9�j؜=�Y��������:����~j_b�7�oj���骔��j��JެWuiLLN��ߵ�E�-�R&�nD���3DG0Rgc�����Am0��r:��&/�p�?���*o�1��a*��v����p���Hͼ�J�hy9l�˿�09�2B8N9�W�/�)�^"���[��'��dٳ�b�! ��|Qjl���8�6o���ɛ��z��$���P���zge��{����|m�QI���t����^�OQ�!zGE��M�ѹ�jշ: +X��@���^�cpu��G_,6\��njٍim�I�d���C�T{����Q���ַG�絲���Р"�J>2T4�9��748�V��2a���K�)8���![cdwM#"�b��+�X�y��z{�R��պ_Q��#N��S�gd=6�܄�޿��Rv/8I� �|�ڟ���5���;�~!������)]S�W3��0���o����6�K��&�ȣ9o�2%�a+-�M�S��|�|;��� �a�Z�s��'~�tz�YrtN0X��Qk���m-��|��X!�_Y�2��1:,9E��B����e�C��Ǯ	�Þ����q^QXZ&3|���Gi̰oY��iw$��C�Ni��%���sO�#Q]՛�h�@��9�0�?�M�U��fv*-�R-�`���^���Ny{�O�uڬ\��O���$����w��}
����Ǟ�rʛ����5�<�!3��5�����c1@�BOZ����uwQ�υH���))��:ܨXmZo���X�0JgY8�>����ϕ}+��Y�2��&4J�sU��B�i�3�~�5��͜H��*�B�	nO�wC<vz�2)����x������T,f%��,�}V��w&Ĭ(����@��ۿl�Ti�d%,֖)�>��5��|�Bi�����ں�ۢM�~�}v�ԉ�����&��h�#���H���Gک	�ǎn�+��G��R�
��d�~5� ��C�N=Z�/�4g���a����T����Wx4՟��;���!W^��Y��?�ċ|�X�b��1��*r͓Ԓq*�HO��f�������9���vM�G�(o���ߧ�z�qJNҞ�@�0G�Ot�P^s���ץo�d��\��.��0��5[����4�-5f��.�7�J�6�E}vX1 ��0�F��U������5��8�m`;��2D�4ە���Gݲ��X�G�q[�SP�5�i�{�X��Q��97N�����)Ƶ�� ��Xj)m�{IX���t��n�9��ٱ��x6��[��K�c������"9!wj�=��A�>�����cW�(�Ԣc����:~�����k��-^��[���d���ci��.S��W@�jO��ۖ���� {%��RO��c~���KS1�s���h��g��� &9��